module gw_gao(
    app_rd_data_valid,
    \app_rd_data[63] ,
    \app_rd_data[62] ,
    \app_rd_data[61] ,
    \app_rd_data[60] ,
    \app_rd_data[59] ,
    \app_rd_data[58] ,
    \app_rd_data[57] ,
    \app_rd_data[56] ,
    \app_rd_data[55] ,
    \app_rd_data[54] ,
    \app_rd_data[53] ,
    \app_rd_data[52] ,
    \app_rd_data[51] ,
    \app_rd_data[50] ,
    \app_rd_data[49] ,
    \app_rd_data[48] ,
    \app_rd_data[47] ,
    \app_rd_data[46] ,
    \app_rd_data[45] ,
    \app_rd_data[44] ,
    \app_rd_data[43] ,
    \app_rd_data[42] ,
    \app_rd_data[41] ,
    \app_rd_data[40] ,
    \app_rd_data[39] ,
    \app_rd_data[38] ,
    \app_rd_data[37] ,
    \app_rd_data[36] ,
    \app_rd_data[35] ,
    \app_rd_data[34] ,
    \app_rd_data[33] ,
    \app_rd_data[32] ,
    \app_rd_data[31] ,
    \app_rd_data[30] ,
    \app_rd_data[29] ,
    \app_rd_data[28] ,
    \app_rd_data[27] ,
    \app_rd_data[26] ,
    \app_rd_data[25] ,
    \app_rd_data[24] ,
    \app_rd_data[23] ,
    \app_rd_data[22] ,
    \app_rd_data[21] ,
    \app_rd_data[20] ,
    \app_rd_data[19] ,
    \app_rd_data[18] ,
    \app_rd_data[17] ,
    \app_rd_data[16] ,
    \app_rd_data[15] ,
    \app_rd_data[14] ,
    \app_rd_data[13] ,
    \app_rd_data[12] ,
    \app_rd_data[11] ,
    \app_rd_data[10] ,
    \app_rd_data[9] ,
    \app_rd_data[8] ,
    \app_rd_data[7] ,
    \app_rd_data[6] ,
    \app_rd_data[5] ,
    \app_rd_data[4] ,
    \app_rd_data[3] ,
    \app_rd_data[2] ,
    \app_rd_data[1] ,
    \app_rd_data[0] ,
    clk_x1,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input app_rd_data_valid;
input \app_rd_data[63] ;
input \app_rd_data[62] ;
input \app_rd_data[61] ;
input \app_rd_data[60] ;
input \app_rd_data[59] ;
input \app_rd_data[58] ;
input \app_rd_data[57] ;
input \app_rd_data[56] ;
input \app_rd_data[55] ;
input \app_rd_data[54] ;
input \app_rd_data[53] ;
input \app_rd_data[52] ;
input \app_rd_data[51] ;
input \app_rd_data[50] ;
input \app_rd_data[49] ;
input \app_rd_data[48] ;
input \app_rd_data[47] ;
input \app_rd_data[46] ;
input \app_rd_data[45] ;
input \app_rd_data[44] ;
input \app_rd_data[43] ;
input \app_rd_data[42] ;
input \app_rd_data[41] ;
input \app_rd_data[40] ;
input \app_rd_data[39] ;
input \app_rd_data[38] ;
input \app_rd_data[37] ;
input \app_rd_data[36] ;
input \app_rd_data[35] ;
input \app_rd_data[34] ;
input \app_rd_data[33] ;
input \app_rd_data[32] ;
input \app_rd_data[31] ;
input \app_rd_data[30] ;
input \app_rd_data[29] ;
input \app_rd_data[28] ;
input \app_rd_data[27] ;
input \app_rd_data[26] ;
input \app_rd_data[25] ;
input \app_rd_data[24] ;
input \app_rd_data[23] ;
input \app_rd_data[22] ;
input \app_rd_data[21] ;
input \app_rd_data[20] ;
input \app_rd_data[19] ;
input \app_rd_data[18] ;
input \app_rd_data[17] ;
input \app_rd_data[16] ;
input \app_rd_data[15] ;
input \app_rd_data[14] ;
input \app_rd_data[13] ;
input \app_rd_data[12] ;
input \app_rd_data[11] ;
input \app_rd_data[10] ;
input \app_rd_data[9] ;
input \app_rd_data[8] ;
input \app_rd_data[7] ;
input \app_rd_data[6] ;
input \app_rd_data[5] ;
input \app_rd_data[4] ;
input \app_rd_data[3] ;
input \app_rd_data[2] ;
input \app_rd_data[1] ;
input \app_rd_data[0] ;
input clk_x1;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire app_rd_data_valid;
wire \app_rd_data[63] ;
wire \app_rd_data[62] ;
wire \app_rd_data[61] ;
wire \app_rd_data[60] ;
wire \app_rd_data[59] ;
wire \app_rd_data[58] ;
wire \app_rd_data[57] ;
wire \app_rd_data[56] ;
wire \app_rd_data[55] ;
wire \app_rd_data[54] ;
wire \app_rd_data[53] ;
wire \app_rd_data[52] ;
wire \app_rd_data[51] ;
wire \app_rd_data[50] ;
wire \app_rd_data[49] ;
wire \app_rd_data[48] ;
wire \app_rd_data[47] ;
wire \app_rd_data[46] ;
wire \app_rd_data[45] ;
wire \app_rd_data[44] ;
wire \app_rd_data[43] ;
wire \app_rd_data[42] ;
wire \app_rd_data[41] ;
wire \app_rd_data[40] ;
wire \app_rd_data[39] ;
wire \app_rd_data[38] ;
wire \app_rd_data[37] ;
wire \app_rd_data[36] ;
wire \app_rd_data[35] ;
wire \app_rd_data[34] ;
wire \app_rd_data[33] ;
wire \app_rd_data[32] ;
wire \app_rd_data[31] ;
wire \app_rd_data[30] ;
wire \app_rd_data[29] ;
wire \app_rd_data[28] ;
wire \app_rd_data[27] ;
wire \app_rd_data[26] ;
wire \app_rd_data[25] ;
wire \app_rd_data[24] ;
wire \app_rd_data[23] ;
wire \app_rd_data[22] ;
wire \app_rd_data[21] ;
wire \app_rd_data[20] ;
wire \app_rd_data[19] ;
wire \app_rd_data[18] ;
wire \app_rd_data[17] ;
wire \app_rd_data[16] ;
wire \app_rd_data[15] ;
wire \app_rd_data[14] ;
wire \app_rd_data[13] ;
wire \app_rd_data[12] ;
wire \app_rd_data[11] ;
wire \app_rd_data[10] ;
wire \app_rd_data[9] ;
wire \app_rd_data[8] ;
wire \app_rd_data[7] ;
wire \app_rd_data[6] ;
wire \app_rd_data[5] ;
wire \app_rd_data[4] ;
wire \app_rd_data[3] ;
wire \app_rd_data[2] ;
wire \app_rd_data[1] ;
wire \app_rd_data[0] ;
wire clk_x1;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;
wire tdo_er2;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(tdo_er2)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i(app_rd_data_valid),
    .data_i({app_rd_data_valid,\app_rd_data[63] ,\app_rd_data[62] ,\app_rd_data[61] ,\app_rd_data[60] ,\app_rd_data[59] ,\app_rd_data[58] ,\app_rd_data[57] ,\app_rd_data[56] ,\app_rd_data[55] ,\app_rd_data[54] ,\app_rd_data[53] ,\app_rd_data[52] ,\app_rd_data[51] ,\app_rd_data[50] ,\app_rd_data[49] ,\app_rd_data[48] ,\app_rd_data[47] ,\app_rd_data[46] ,\app_rd_data[45] ,\app_rd_data[44] ,\app_rd_data[43] ,\app_rd_data[42] ,\app_rd_data[41] ,\app_rd_data[40] ,\app_rd_data[39] ,\app_rd_data[38] ,\app_rd_data[37] ,\app_rd_data[36] ,\app_rd_data[35] ,\app_rd_data[34] ,\app_rd_data[33] ,\app_rd_data[32] ,\app_rd_data[31] ,\app_rd_data[30] ,\app_rd_data[29] ,\app_rd_data[28] ,\app_rd_data[27] ,\app_rd_data[26] ,\app_rd_data[25] ,\app_rd_data[24] ,\app_rd_data[23] ,\app_rd_data[22] ,\app_rd_data[21] ,\app_rd_data[20] ,\app_rd_data[19] ,\app_rd_data[18] ,\app_rd_data[17] ,\app_rd_data[16] ,\app_rd_data[15] ,\app_rd_data[14] ,\app_rd_data[13] ,\app_rd_data[12] ,\app_rd_data[11] ,\app_rd_data[10] ,\app_rd_data[9] ,\app_rd_data[8] ,\app_rd_data[7] ,\app_rd_data[6] ,\app_rd_data[5] ,\app_rd_data[4] ,\app_rd_data[3] ,\app_rd_data[2] ,\app_rd_data[1] ,\app_rd_data[0] }),
    .clk_i(clk_x1)
);

endmodule
//
// Written by Synplify Pro 
// Product Version "Q-2020.03G-Beta1"
// Program "Synplify Pro", Mapper "mapgw, Build 1618R"
// Tue May 26 09:44:56 2020
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\e:\gowin\gowin_v1.9.5.02beta\synplifypro\lib\generic\gw2a.v "
// file 1 "\e:\gowin\gowin_v1.9.5.02beta\synplifypro\lib\vlog\hypermods.v "
// file 2 "\e:\gowin\gowin_v1.9.5.02beta\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\e:\gowin\gowin_v1.9.5.02beta\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\e:\gowin\gowin_v1.9.5.02beta\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\f:\gwip_test\refdesign_sdc\ddr_psram_refdesign\new_ref_design_v1_9_5_02\gowin_ddr3_memory_interface_refdesign\ddr3_mc_phy_1vs2_2a55k\project\temp\gao\ao_control\gw_con_parameter.v "
// file 6 "\f:\gwip_test\refdesign_sdc\ddr_psram_refdesign\new_ref_design_v1_9_5_02\gowin_ddr3_memory_interface_refdesign\ddr3_mc_phy_1vs2_2a55k\project\temp\gao\ao_control\gw_con_top_define.v "
// file 7 "\e:\gowin\gowin_v1.9.5.02beta\ide\data\ipcores\gao\gw_con\gw_con_top.v "
// file 8 "\e:\gowin\gowin_v1.9.5.02beta\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
nGQjNTRggZWOT6sWc6oyraDUFLfWAO/HbLF6wXbCqXPNp9WCDJpv1rHVczOIVgncR/b0+UeSwebZ
OxlPzCeuO1qPl8FPTKiUyycPd+J0aSTr5vl+//g43DlAnrAZWpp+9NwkyX7Tl4KQV38q+/ZFnqAd
fKrxDpwkhDu4v9GmdKTtVryneeZJtk+qfqQLeux8ui4DI7WokBCiLCcnunBZc7zPDJ4RNHhhj/d6
kphLiA+2e7BZhQi3+S17OFvZZeAZqB9QHyWn8tsgCw/p96pTPtatJ/h1TGMYgxgbBmCeWweLMmye
bCwg5pbhghYptD2zVIQFJWuiylXMfypQ3ZpFdA==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
x5gHfLwQ9h6IkqXYFQsKYOoMTbgAOviKZwc0Vf339pYT772gCzJCT3UDF+YsUsYbK+Pq7BKRT6Uf
HBulNYuf7y+Ku9k8h5gb4vT0dUa4DG8OSdHb7R0AC/h0AeBTlns2hBJ4OSQGxyyNBp2s9HonSdOM
8ZWZFAphVVtPxikUpfU8q9qzyHTb9jMLF3VfqHt1hy3qcsmu5t+UPmv9c2zjTl4NXRMUl5483dXo
fMq4baFS/ju/wiHFuRhteazMg0mM6BfGhtM2aDlFaVzlnFbwItgar6Mu4Fk1u80ynR+wqXfj4ur2
96zU62Pm3UBbG8dYUGOAgfAhYDkhAs6USGbytQ==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7104)
`pragma protect data_block
bHbm8M4o9I3o/LZ6Qfxvvulb8QFxs1VkIzi11TVjvV0FewNSw4catw5WtNyUk7HamThcQyRqr+YN
pBFi8MZQYHezYX3inYaZ6h8JyxeLlojBmH33/e9YOcsTdYR3Zz4b49M/cDCPGlsTVdLKCYcl2g5Y
oIIe46zzx48pW6tIYJ2U45EXloz5ZTLseu5SL5++mRpwsmDEYs5hPkimYCzBMYaw8VcD/Z6aC3Mi
3UIPxDQSB64MZhT/rkCi2UrQTA2ERQ9hAFjlSeykHFO1/MmhJuZLl8K0vP5Z4//9hhxJzu3nCVsE
xEfngxiZs1RrC9ehUO4Z6Gk1KUz80k0O26dO4JGkEMsrxv1idfTvI3VX5NDz1r74PpuBUY+psKGp
1rs1AiYLzrYypOYnul3oJEduI2ZHPmTg5alRWKR7qiIJ1vqWLJl9lclGscoJRY6SE5d61nGha4lx
JnIQORw//8gOVRK164GuD8aSnx5+YjVnTtdBvzLejA9A39JfjX8BDfoVi6xf+LO8bPbXzg4Gog3Z
1lyewhERTYEeh61YoLIGDdMjOMsbxqNX7ThgmHvJQnoDqscKBpNjLGMraqNiP1dzCi+aFJXIZ+xc
3PfEO0C/HqH+QWJ/LMFT9xmRF3D0uCe/hsFK8BC369uXagceLNsSYNjmzS4bUsmmExF2+RIuB9QL
FjbVzegdciZnoUGZSvx+UnVjtN5HJCdZ6XOsnui+MekIMXjPfzQb5k3oiKy2L4g1+OKRs3rL3nG5
yx1MhK9vdWCKUIR9QI7HDrCfgMZvC0L0WYABm6tkYiwCgUAv9zVFHTPFbCPnWF2ummFotfr6nZym
gu5Pp9LUUBshAaZHar46K9OxYnj2N+7zvw2GEGbsS2Rj3mQhCVI6fbovWZornCj4IzCdTXcsFQic
xRfjaHB0l6M28AH4865dJfpL43wMpXMBZBz3K/ikohZ5QhZtIk5F1Qg2o1HtOZqGrQTPcj0Gq9tr
ftJWWWqR+2Hkafur5md/W7jY7fU26+cTOVZH5z2C0Y67PcYiHgogMObrNcSyI2JRko6fEkmG7Nqt
QHbB/Tjoea0CQ+WJdoKKNbvwByZB89TEsKibFFaEk1axrVsQoZ2TKdJ9d4Y2COJVFrUbM+8eCGBW
VpsTxtzWU/X7Rh50h/X4TJhS1IFrTpS3viI+Dfq85iUDgc7E+zUxURUWA3nZNDbdRtU6GtdwRYzW
1z6SyA/RmoU01H7fdygQPKNnbAGXa+zM+IINy2Hl4omvrqz2Tc51bHmJx4+FF1fvsNRIuGWYLcXd
alnWEv6BDwLxeCRq6m5x+P27kC+3eIE78PshHbliD0QktnNjEvrmlLvxoutX9U1YeSCyFa1by15T
rEqbSpLagXhQ5ZIG0579aESOaz2T8E0IULrX0idyGFjIgKMWc3uj1aV4ux3hpQ6UqPD6ZVUaqnt7
3nlgS+IbfCQnVSfV2yvTwSze1XaWUDLnRyC/xCZRdi6nJw6Gdcp+fX9ngyYx4ezQTgW0L8/kos5c
lUhmD3nCyhh+95QGJodCiS24NJtWQ+rQaWX5nyz8gv88561ZcxNUJLu/GvkNbTNaJIlrCbAZX8kD
Fe6q/XYb30m0MhsAhRk819N/NyQUVE7GrZvWZGv+sKJgI+72WNoeHOWcDf+MjmxKMsprk/9Nornm
LLdsA5bqb91kUDQGdwRCTkjuYhkCNDsfrJ1gbxhqW86K9I7ZTmIjN8Qw44LphqvgGCjmwJUw6S+E
s9JKQnzQU4WByr5Tftzl8xDNwPv1rq2E+h6jQCLx7MrYVd83FkguSyKW0xWs1l/0BdNuQfZgshna
pouDbUr9TK9vnxtD4qL18HioAhIKmS1yyUHPql2BJmi3vWPu0zFeQo1XTeME+ebcYEyirzgvh/aE
aTpg9udOQl7Lht5EFgCxx4Vb0gI1tpyedHI+NawxkIfGCa++tp+ZEDLiIou8iZunTHz4wfcxvRhm
S6a9ZpkWy+G6U8IW6AG63Dq4nUr+iwqF+GeWuMVjKUSGgh7y91dUekSfF7n5XmS1TLeRRvPp5obf
+09izZmMkWO/2DxayZS2aDbFsiFObyQFmE+fk9zh6sYR9F46ejNgGdlCpEz4OHj62zbRQocF/fOl
wQDxIFexLJicUbKOWw8UfGEFzIF5RBbcF6sfOqu9gt4Dp5f7PDNLscpPTUj/+84XTkeUKoYz4HPF
nZScwWgRUWhkK2yQDE9dTa02zQecu6w/O7GAPxvh/ANiIpxCtRh6ig7kXIk7p6DMWcBSGgbZRPRM
UdRYoiuqO6u1S0Z1Qdc2xrg3gNVPQGpxHipDXUDqBA3NbQ+fWPM/woA8zbGV2xZ5DgnV4KiYKiN+
7PZsjUVYI6TX7CwKcN8s5RbvsJk3JUiDe2mGqjX7WiuvyXgGMqAGIMcs74Yymo6/VSYMOlHnXfb2
c5bMOH2IJ+6JWyN/1M5w7bkuWEvY0EcJw0x8ODQz8t424Y29NXXZN+v77bULpVyy4pD14gV4KiWv
Ny+FwPfdMXdZo2BFsP4kWJVDc/7StpCa2vKsHyRTYrNzI6wkd1cwlH3SEQngEr6tqG3RlnZSmeSs
apSVQjL3U5IpBZrUTsdDoQGIqlXllnWe+4Tyh6usEqI+nPJEBwM5G8LlIGPQIKCU2EZ1fpsK0bUn
R8tL0lCmEIQvOPHx7TCIxhUXLdPL0khW1cWT8qlKwoCSMEGsvI36inE4X6skltwDT+hklalnoUry
IPdIRW4/Sxnqbe//rqyCsR8eQcsSPJsmodfdj1h6gZ8TrknvG7VWo7KRUoleyqSQ3XR/lh0ahUpC
V5x0ifeIQv0QvEOMyHf31wTxL9MsXuXj3bW03Vpc+sNstVsN5gZuUUbSG1/IcBYwP3cmt2U00flB
uc4/BG8GuhYTImI00SoLfHnE9i8OKIzcEC+8a82A9KAUPo9ggFubX3ZDPgqswN6YVoXN1UMtVVSP
gLkUR4zD+PXWUZrvQA9kHvaMI1uD8iJur/3O705K6hz2V0tmK8C16SStKI+FO8jgMTtNIR+PdvSf
0EtDwqlmht05Bn1PmNATujZd3TMvT8xV7bneeJ5u+3AZansinNh3X5IKVRyze4VvJ1i+4vK0wblV
F0xi8C9DvUUqBgebWByNvp6TWWwF62px8ATCav8HRyfRYztnGSj7yfvDKchby8RYWqmLir3lAE86
BChQMmdU78cYn21h/I3c3T7x4C3+kKccNi/t0h+VG6RKpBM9xDvCEuT/dvS0aRCp/tVdPIKIAxuX
v22MIjXWV1uWE/dWvAF6qM7aUcjb/UOokUupoDPimY4UMX1AUiNugq2EZY2zRKyleKnlznbYI/CY
RSMwuUkRDX69g2Dg6YuoyXbWWeoND77XjN94na2qbx73cB4gpDovuZopzaAq+f5XGMM7gwDAKp5D
pATlaJei6znc7UXqfjP55wel+tGc/viq/agazF4UROzu2znQf7rEH6JWR/Nv2V/L/7TqAhiEvZvW
SGcBIBbOSLp2TKQARL5Mtem5kktl44Xa6US1yC0eMN3Ee1TCeuwlmy67/6VdEN0VAFcb0+iyNt4y
nw84b9NvlZc5i6lkLVo82WMrlp8ibhgm+PF8LWwPmBODeM3Atgk4UuYRPRpoSVXR259mwHqXrNCm
6bEsvZIHT7lSDtRyf7fwVkdc3GYONH61YxVW6qiCNyZ4+QkX7HPGCL0qcFS9+5e1fvyxChAlnVbs
fGkLZ550YZ9deQrRYbogXDR4OSidWHDPyRPbMYjBx1r6Wdps6BE+3rzgGZ8gk82vnsrLcX9bewtG
RBnrAm2FAY22wAZTNO/zRbINSmYMWo23NbgLiZYNw+lX4ATW4svuDgq1DM0+0pHAdFcmO3IuXtfF
QkPc2PbvVdg2bvaKuCrbkVwcrjZjLsSTmZcvIL3cZosAJXyfRva+8QgZ+x6hJhsfX6Aer9AcBWN0
NvKqFHjAwpMCmTuzR+mIzRCay4eknmbRVhdEol6hRiigtCeE4hAjYwsQMwtLih7dKYA6gUv0PPGx
gHwYcCgJmLnH7gvz9VKJPHBr9vjgOsI3FkT1MHgCMhBoJKY8a9foBvT32I8XyCA461zUm6+2+d5e
v9OjxXWnJkLOJo4s4VDxxleptcs6yjXJr7QKO88K87H5855okjjhi5tyOpS8gxfx8KmNXrlZzokK
pH3SUUMRyzLu6nJJQnd/ifuXCWkXL4IR5+Cs1QDC4y33SSwm9oF50iz7qLkTMkwbw7+lmCzWLCb6
2t+LtwLTHXecvgN34v4gG6kAvMLjbk4CPppksIC4nXSaHGVG+R9QnAxUaWAVtS61tl2G/w4hjmvU
2UjRrmuK5w+AC8lpas2cqBVwRIQ7Zx5cg5MFhiQMl45pWOerTRwQzMUoY2fRDRsxmSpAEhBIY+RJ
SCJB/H9Vj7P3hceZ7huidD5AZANYIGKLxtnpos+451q6baBZVK2HcU5w6i9iYhogso/CCNvdvEkK
3pXMavGiTKzTpCUUl06y1lfvOLefljGDPH543E3P3mtkxV+zAe8oYcF34BS8/PzY/sa1w1jxwp82
VQL9pxy0taGw1BkgjziXx3sfGB/l3ISESh6pRG8Y26fYbzJKOLlGsRilwWh1z7ATJaJgTI3AsX7J
flQEc0r1NHbxZzgNfuewwbWkA+Lud0qhrUxVE7Kh2ACYuATZQdviCRCVy3ZGezXYWfG48pDNG5BC
0vHByIsGWr2IJF6b9GwHqwBLsBiQSCFPU4+Xbq4omcSqwmkH1z8Vnd1Rv9Z2XWH/joHBs4+ASaQY
MP48gXFcf2HitT8Oo6CJegs4xwHCRQ15VKyEn8xSuB6nJUUNKbiNnndsT/LL2NDC1h4Kp7ecXEIV
6jmlNy5IKSHzMeGfhAgep0sEeprsIGBDI4qgPheSFW5RErE5u8moLXLKPumUxtAIQF16Yp+0IKbJ
VIKmAO9VahJ8kmghlhHuwxbiJdGAQp6gdGPp3tcSQ5e5P+8qbiUktX2AZqhj2KWIHC6BcElS4UXL
TWq9DIVHQhf/ep09yiHyBRLXYgcWL9ATs/8GVCeME6uBm1PPNsBREzkURYJ/PLD88YI0bVX1QKu0
TLdCSEmmt1VGwaE9QDyW/iIas7zg0MIVK3W4aYEWHiDF8yufHOtB7lYcKGn/SnB+81xbqfTdRjd2
8SGnArPqkE+bMNS2iM4DPiehj13oo2253rL5RI27r5Im6CHy/EwaCgOILA1q8uakDxSDu0O3A6Ca
8zmWlR9pufiaqclYuij893RYeF4+dRZPelSPi8lGtGsknVh6kyHBU5Qbo7td3w7OMvDHX2MJceQM
0qVo/jGayQ90rQ+If62jjLYDVcW8AQHIpQotQpiK9KAnXvXiuttwyJoZixuCjvL/fMEGQUR7NPij
IDhI0VwpCQIqjar3T490GQrT+P3fSxzuoGAfOdGh6yPEQ1ixQPq4wk1LCpuuQLwk794MrJsDblf7
wusLrBc3d87IVCwUf4oESwOcUka7Co7Uf+RmdGstBOYa9T+Ifk6xPYMIDNwDfEft07dD1tB2ylNn
U5JlX/4LpDjuMGqxXCtz/UG5ww7xNf2Jydg4luGraaa2ly7RBeOFqJ2f6t2dSMcFvYYyrrSZL/Ii
GyspdN9nulqBtrOOUW4Gc8waX1gMAVyBE/E4l8pM6201ZiWDP+RmJtg0O+wBnpxzlupHtIn28HdB
8CJ7llxfriijkKicR8e6D+WC0oc3xYVMfGA1LC1ob56coTOdYqyjLdibeHxGs18F2dlmtX5d3oMC
zUcvnCtU6ocwDHiihg3RK6YbMsbYj22Tf1/+VEmz2NiHTb8maYDqGBlIYlflbVcm9YWE+pclpURv
I9ZqEmK6T8fiFsCMSY6ZIDeTBFG8E9GSj5azvIP+gqXmhJ+6yXrYBFjIMcm5TnmCjI0JXycfvoub
1IFN429Z/vGT+mZl/JosBL+kHrHdz4Uu3QrzQ4BNhaEZq2/n5Ytz8zvQLReSalKUBBITm7kT/oUC
hq26tnfpNfgzEUDYdp4sMq+JZhjw8QMFgJ5hw5INsHsO3MIy5tp9jxguxwzRIE5q79p9OJ8GH4Oz
PR7mA6x8aMqeHobQSb5qL32gACnTRGaZuAr84ignqh+K9/3xC8dpJsiXzsREHLSw/vp16lwaFhZ/
fT6ZJyt+I0BxcOZHtnJ7Nl8n5wVhrOrBbxYG/OsAKbOwtky7erQqi82SdBZPCu23zqGMoGscKZac
2ZFI6/K9OSwXSEB1qGfxTAGta8dyHCtGTvq6OcwXgdydCNHvAjq85zCXoCWZUdHFdvkQAhTNqs7B
4D8eZODvXSUS9CgbJRRB0zDlfaqI5QVHjYv/zEGdJK2P5o1MVLxi2J+4hLSwQ+niC5I2vTnfo0w/
6rLMakS5hSCmF278qS5qVRRin1tYg6vq0e9hyhCGWCpNOfL9ki5u6rJ213cnTSrY0RVV0FnaPYcS
7huXiUpjDRLreltZpzh97nLBbRrbuxulHKXzBgT0HFuKgiCu3o3oC2bSAeyLhHHOCPaWE14jbzvB
1TTzkTNl21MoMKClv1W174/xsqYV8Y3SkQi5QfOLY7I8qaF0Jxea1vNfhtoNH4tYiKAGFzvslh3T
mH2VRbcCxI1LNJWhB5tdMGPo3zkVHNLg0n8oF5feDN6CPkGHSgLN5HzqYopEjrgnbODRrm4X4aUb
k/2m+hchm7Mx/lSeb/CfT5vUskDxGxWBfZtpxGpGarDds/SSFyjqlks+xC3Dnp58SJmw2pL1AVTr
ZNKQqe5K71nUoTkO1daiJh7Y6mbexSAU7JUKVX/E+CydyF7uBOKhkSrbLIzKQYGAi12K5lco8Bxv
IbAP0RRqQ0mxNaj0gsWJoFVE/bI/VSdgIEGLNcL4wXtqmt8IBsk44dOB4UjuFqHQNVfB9j7kYpiE
bE5quf+B7KZT8MbgZ9oaxs13xIS3pegmmTKfy/cYfawM1dmcrIXIr3wddvvUkikzBJamEJq74Si1
sNkfF9hdippAQKHHhEju/uLcmvlDJDbTSmr3Dqc8rmvW7M7RMvmWQJtr67d96pcLtqouY8f6Qsfz
U5lsJTlZkcg5fvHqqqq8oBDjd91s2psr8/JYKIJXQMfpjKOhdAtSVicCv2xkJ2IZLMuq7Z6MsN9Q
z82TB/DS1AcV14whgaixAd/TqLX9wJIIsIqqHvCYrNawGKbm38f3qlYHzx7aSJ4/B8f7ujGwa9Ol
iXFRRXQInhjCrH5b2ZWOYOw5VDAR6GQTHKOo0PJyyy9gWpucIDgJg16iQjQLzKsjBjmeUGgbp6mz
6bZ8k92cc/n8H3jjxWbzXwsHJBzkfJbNHxMpPHylwikFIft4BD3wKAF3RkCn1JUSSnbBOqO6nGtn
/M0x6uucimDpIBtkpi9YKSix1YT1mIdUD3nd24rH4eUka6DRTJvxz0zFmSXr621SKMC/cPi0J8C/
Te/4e3eHXMawQElCoSY4ZXOPlsV8cSFuJH1YXvNmA8448RIbg5ajBKLetNvDpbzOB08tKEW3ARcT
HIGY8Vl8WgVWjTtVhowrPWJf0yE7MllO1YgUddZRO2mL6DIXzRR2ltbJkBO2Eo5NOrqf7raA6ltl
4Aq04tlP35j1j14V4Jie+RsqjBLJrwmO82PTsuNSs7CUeIVQ9PIiGOTkPqCz7S71xh5Xe4fcnBKz
652W3ytsjVSUhmNPanOJ97Mn4K0B3KwMFfYGJRRxaLKUWUYNo9O9/re9eQ7VLqXAmW/t8rx5peDk
mJFsj0dQpU1F/IXM28ki52GIIEzwlNHvbPYCGlLuGypXZj4wO8C0YK1YqukZy7b89ByAJwSfR0mv
IJH7/eeJ4d9AprW8hUbh+Qkjaj1FtS/nszW0WN6gjmcQSwGTCD513BEwXQSlDmIAEaV/rdJaTbqx
Cg2GSDL/Hlmk7iAEiZ++ZT3MFaxjD0KT6IjDX6KRDVkOmDKy6b8Iui71IbRP0fNNcjq+n8gmXpLY
8oOQi3KU+dighO9OsKyUK3d8yFxA+DnGyvlrvD0ldgdwoMPSev1uUW8gOhvXsnGJopW//SRKDuva
8tEQ2oijK+DDyoIDEn51UR5Ji8F2zyNNAZhv0Da1Gc8jEbU147wImql0wZW/9WSmkJBnZE9w48P7
dbutg4XJigtpfaxudXUmIb9Bo+VXwvJMYxxngGo+xBTBC7SVFvI8rSRRL57/r5xDJhnwIIivCKsZ
0uu297ZfYLxjIGrkviajJIrFIuE34SqDlLepqUG8IeJg9k4ZsoVUeLXhTjMJx5XgsZBiZ0GTmcoR
0/0gmCEASouvj2Gu/dIfHp7KzjOSPUNItUiqAV0A5MjfLJ/36xvPRaB/ngaSGqblncLEApa4+HXA
/SUKLzKssJgzen/eYEeyElutvb+5wDO9q+kheoL/fkw2B7W9ec9XLJoG/rRKHMM3nd0EiTxUPUKq
HQRZmk1y49vbOZNt4RJkDdYjTkV0LQQ5N5PP6QISGJzwYeb9LBCfznVVciCutI65sUgFzZhcgHLk
52E7wE3+TmByUP6K4oBff0kUIA6E2ITNkx7Qv1QJ4GsvuP4Yk6xP2DBlWNWqQze8lhoRUlrVsrz/
tUtH/GBa1oGPvb2SzlrgaI7tB1OpurvD6vy/KnItajkH1mMjr26g1SDfAqRGUUsipj3H54kXdF46
qjp1KgGJoJHN17W1KSotzx3phZ4uGddZVQ3j5CD2GIHG9AYY2TTEvSNG6ezz5/MpSXCLTjc28TRh
i/pH8l8hswnFkM7+PNiP/hkKMtrA6oAcVhPdOQt7GZoMoJ0iL9KzeD4YJITKvv4CI/6QQ85rTIbp
WhOSFu7NLzSemZSwNV9ZEfmlXiEDEt6C8fb6qRBTzE1w0HiTCZUpAmDCS5ralb9ZXpIStccseSgW
JN8W0LGIXHiC+ZeXBuPeUI45sqfpXZEJYvkGxaLfRBEx++OSxDSmOTP/349bXHji7BWXJuSnrqhT
/lvQqY5i5lJb1miLUTZqXBi0zUvMPbheOBULWlCkRAgd+qRUv7v6ZaD4bVrpXCVpQ+S1cKIGq671
KUinN3pwh/cxCuDkgU7RhNvjPI83V/5u5hjSpJ7NHNEGyDDeq9OeClw7TMDPAPG8zMLiJUqd1aDv
RphQcLE39wGCptugys8lCMb7i79z5LbfvhN7QbgAiwZnGxW4wOWnVDrLtQjZmJXp8Wnp3Zs0/4p9
V4V3gVSWL/CcQ4MO2OqmfwAHw3K6WLIr5tJVmGKvO/W0qyPI7IEfeuwMCuRdglaTqZ2fDMcrRDfk
xj3A5n/qDRwdvpEKfaYYer/HUuNqXKBaNnKdZP6/XsBwvETIpgE1ENHbjQunr87g+pMCHygvWWpO
z9zTFfJ3TldtbGOL+BO3LAode3bhx8o2F2PVtRW907eQ0JBL0pbaX0BQ2beyML0QctakmRewFT0V
iBzlCY6RJGMNFzubscbc1Z/b4lu36Zi1mAeftbbeiqQ205U/
`pragma protect end_protected
//
// Written by Synplify Pro 
// Product Version "Q-2020.03G-Beta1"
// Program "Synplify Pro", Mapper "mapgw, Build 1618R"
// Tue May 26 09:45:24 2020
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\e:\gowin\gowin_v1.9.5.02beta\synplifypro\lib\generic\gw2a.v "
// file 1 "\e:\gowin\gowin_v1.9.5.02beta\synplifypro\lib\vlog\hypermods.v "
// file 2 "\e:\gowin\gowin_v1.9.5.02beta\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\e:\gowin\gowin_v1.9.5.02beta\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\e:\gowin\gowin_v1.9.5.02beta\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\f:\gwip_test\refdesign_sdc\ddr_psram_refdesign\new_ref_design_v1_9_5_02\gowin_ddr3_memory_interface_refdesign\ddr3_mc_phy_1vs2_2a55k\project\temp\gao\ao_0\gw_ao_parameter.v "
// file 6 "\f:\gwip_test\refdesign_sdc\ddr_psram_refdesign\new_ref_design_v1_9_5_02\gowin_ddr3_memory_interface_refdesign\ddr3_mc_phy_1vs2_2a55k\project\temp\gao\ao_0\gw_ao_top_define.v "
// file 7 "\f:\gwip_test\refdesign_sdc\ddr_psram_refdesign\new_ref_design_v1_9_5_02\gowin_ddr3_memory_interface_refdesign\ddr3_mc_phy_1vs2_2a55k\project\temp\gao\ao_0\gw_ao_expression.v "
// file 8 "\e:\gowin\gowin_v1.9.5.02beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_crc32.v "
// file 9 "\e:\gowin\gowin_v1.9.5.02beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_define.v "
// file 10 "\e:\gowin\gowin_v1.9.5.02beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_match.v "
// file 11 "\e:\gowin\gowin_v1.9.5.02beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_mem_ctrl.v "
// file 12 "\e:\gowin\gowin_v1.9.5.02beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_top.v "
// file 13 "\e:\gowin\gowin_v1.9.5.02beta\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
DI4rXVSqQQakdxUiFbNMpUcFqLtxiH/v9VC2fotO6RT5oJx4ujfd+d8ntglwi9SznfUhuCDdANfH
XYMgV7tqilOQ2ZawjyjFzCrZ5SPXrGgsruT0nRljnPbi6qkiFtugOcQTRLawx9T7//cBM+KloXTA
NW5UEesUVY6XIevfIUZGJ1ure5Ny3juAG8DwrfgVKoVsVbpFHGqkn14/CuCrPfgd3cNIeMnz2tdU
fIIQcJuw7/y7oxsPIHnSNjduB2VlABUbTul3/U+MLlIz6QrQXnGGd0gsk0VzmjNw5t92AUKNXFJQ
KgZfLCLpjgQ/ZbGsMSNTxIFdLQdlxHMJmC0vaQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
BJq830S/kOcQBA2JJ2q4S6I8jB9jjQ+2w4M1vD4Tqw23sKPDOhifxjr0/o3W8kskkjrPH5ExmJnx
4+Ax8NsC3/y94RfnMYtaR48dVDd/uZPC+H97z8xQbMlRtAPIPBxmvbm2XF9esKwvNQk33qXslMT6
Af5S+VRtkbzP466p8XNJQwyztsU9oaM7FXV1jV3HosbJuRzcKVPEOmo4Dn/DOSxaP8rd5LPjoLqS
+itgiiOB0/sBM3oF4lMqNh90Lt7h7dN75Xc5z0AOiCtIi7ReGbnoPIxpLrTX3YY2f7/TaNJjwe2m
A2muDv33kmPJYj0Qn1mVE7WUxAUWY5au4KLJvA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7568)
`pragma protect data_block
8x+JNuZx88Q20DctkrO9OTxw6UVUAd4wY4s6SbOwa9t2nOHXdHwsnOAPaBwv/kAA4pHfsgjunsZR
O/IQGpkZAQrZhUFGy7uEaE0o25Kh8kMyNGoKrQ172uQSH7Ml788IHbIthQ7F6wvrVp1ZC5a0FK1E
DMP6+qPvfHCyjn/yBMSJLcuf4I34me05TbK9hHrypOD2gar7+jAkKfurjvhdr4EgGvnu0pnRB4mN
sTS71HsBW7HpXTiXEmwC6DwYwJtviKwk0rWSm+sGldkAsnxcye0iWcnEpDykgGjHpzCkzIMu0RlA
BOnYabXXbT17znti7KOt23dBA6Ms4tLNH6UwWVhOBUEehXKeStkFKvbJOP2Imi1V/D/iZArBcjcz
ZjekNygrrcoK6Knc4ugegnTkTEHP9wFcfaCM/0QPSQsXKpI3djvxipPfEc9y2/hfN5twZdN2tkWS
wWtdcGY99N484CO3u80FI/23Ql9DhiPGcPQWxgacRL/5roKvG8CQxv+UCLEUBdCjQ4zggat93DVg
mcvF50T6vMRObdY0HPZuiFUB5cutuaUCkW+ilttL8BUhy+COdblBPwbMODHmt26XY6ucNP756Oqc
m00hBlAiW7/L0whjcchxrGVlVDwARDFHd0k8I1p5BK76BKEVu1pOMsJBFroiNkXtubgsGwNH6kDf
4jrjIf+2Ucw4GrrTPmhEr3l1ipFU+XSBw2b1ev6qT7HTnfk8WfaiIEmcuW5iF950zOMnaxcvtBhG
JTM0bKEFw1s6ikljxO+T/n0N0bEr1fOIut7PKZJou9xa7YXgB+qpxVrPxmTQtFWtEzBoG1kcCKJM
B9uzfJmGXTjq2EC0CyyGCqncsozKs1dvhHGyFY3rKd0ZUOU/YA1TAWxZWQL7k5P5ha/hKTESn0/3
7qpory9sob9+Gn3ovn2R/0nhHrLO+t/LmkLjttNG4gWfD4Wde8f7zvVtkoUi6teiDWR2FPlorlrn
kqp+m1Mbmijz4gen4ezHXFDsohzBzylJj0Ytrc/JRIkJYHvKhfIZHNOSA/VOD36iCUAoBxgC7Tmx
bdOsZwedBDLEE3SaX4rlTN58Myt1NR/UXFLM6XtxFI10GuVfwnnTDlGg9d65eSwP5o0vb6AUPmLe
iTAVVV8xXPqBIW4paIrKV6m4oCwHpsn0AvyQALDPoJRToeuEgismACJE0wBjVTCqByUF7tXTW3cf
/ioY+rRlX/Yo1+K7NTmuANLP+TEP3lwe8Kfysb84ghNRfUx5ktxPS5GCC46JRdwclfQTiypbXNKF
LBMokUPCyKnwnVFHq/8Zb6h7tLQQcpoLRkSNhies+bYiMoVvVk6Y/4qYBK2YaxWoYDZLu0OMtU6e
lcBLxCK9AFt7cvVDMpkxsTwsN4bB49aLpOYp0c3lDGVL0b0l3OHR8kYBLe3CvstzSOssuoU5e/NE
zRwicyJis141vWe18nwJ7XMUI1p+B8zHe2E2l6G5FPTfOegIMLlxHKmSaCKegb0CmEIeFyi9t6Dm
/ppFxT1V9ztUcU70frSHAL57zgMTXHB91pgBIJ0F4RrrBrXhVEM19P3cayKhbDoXwXcEGw0OSa24
pTBEHmI2/1sZuM+kpYX35B6d7pEpGeVRSOtG/PAr4nb6qxp1l+OnydHD3Jhd2PyR7wPeZ9VFSwgC
RNSa+YQ3XhLGnK5Ep6j78qhGS8YAVDgiyiJMvSYns07Mpy7EIp6xtR2Tzyi/IZ90KfrRDFwjkXog
KCBIhCV74odUvNPEqaSX6hOANm9QlKDrMKslqrx8hUS0xiH4QV9X5Y/Eyb1Qe5dJNtjASkhihuEM
+M4EemhXEw/YxMkDNoirymsBfoRHXK39AfUPwTmAIqu/39v26Aq5jnkIjPPrwgO0me5pPV0mocpZ
QyEVSfUxf66BR9UswsZmegnjjs5sUB3jZypRWwxFuj9/eOgn0CCSV5q5qi88Ue+4zEV8PSujEjFI
sjkuVy+dWEAihOFNg9QuDDDJjMc7pji/L+HEVT3L4gmNIr29Umv8emMVlkX8OUzDDFa1YNnIfq84
NqYLfPFq8mkH0a47Wp3wpicPTPE+CKnp7Kg0ur1/LlWYEfVuFmfjWq9X3qFa7hRl1z6/n/8iF/1D
t/r+dYiovPa6r0AWbIZ/MA+KokZAJCd1OHV/hyV2kDjsuSkWFssZ/C7468rCIFNI5Stam0XPw41e
AIe1uBWJF1pXfLKdJZ3S5mGMXcKRTBzBV/ELUjs0QUZPKLPuh5YEj5NGAN2TWXcZv8fzQRY1XHzm
DTBcol1q3auYhMR/JJMyHuUa6VC7VGx6XLSCpzLkOlgPFONyFzb/9Y6swik8Xf8HhhrBTPv4DOqm
1G0hEEv0lfiFjadF7Y8vdFwCkaW/JQ8qsotY86WhsKqQ0UfMmx+H10qeZpoio5KFf1P3DbCF1S2o
lKRVG5OBZUrvhvuID1gqwdwWHfx8QFYMAKfsY9rOhJDhoo9TcqqTj57ZLXmClK/zBaU3OZM4eO9u
aWaCziCqE6M0E7wGglOIuIgjmUbf/malD5pBywaygyREcL47ZN8Zgy6ZEzN1SI/vppzVIA+8DjSr
ZR8AhuKBACY7V0W8llk2wIi2IwoUWr3ZEpC6RG6MJtrgvAYUYFkHEhcSKKM/3cSO73AkJ8zlxJnO
E/jQBiRkHND1EScaQvfkDXx+hBf2d9YwKYX513LXsrb5MLpL79XXI9VMsE6A9ygSr9IijHUNHxcC
xcQpXEERUPsHuiI2iHt1PSp1cfldJ0CWPh4dCImdOtq1RW5LorNEPaCu9XGaWSr/8dO3AdLrY6OU
qxL5PDkK/qK3wsDCarocsDwQ1uftneFNc7ztbKPMuKvcf6UBocBO7A6Xf1XHLUAjs27WB3p3XZ6t
MQF4XeakoHRxO8bH1BlcR6QL3uLzH1Arj/IlEFhVefCIrEfCe1vkVPk13y0XblcYb1dvwsoamXDw
8HfEwg161cSzuE6b/ZMouFmNRbvWycSu0/FOGa5/X+xHYYvGSDH6wiLbX01JtXkpasAVQkfyhGSv
8Kt3GPjGMWZj1z/eZnuxNH1KVkTTIUIg7R45YHUhh/GJjnKtr/A79NV3pcKF6qYZpXuJ3KTv6+ly
psk37F1u7Ecuh9GJDCuWkfoivoLnAwYyVus20mSZec8Ovx6sFlh3Ku/xy0lkatPkYa7zBETDSgLm
fPAuUVL2WCamiR5vTSi2Qbzhv4RuAAnHAMmH0TmtBsuzIMTtlk6v/2bVSrUcqSYqPoYDfURiRZUN
sUGeENrBNNT2AiW3n3fqPfID+n3WIBe6jWtihkvwhZ/19Qdf1R/n8OXr9cjlRQN2t3oZP9tP/hsP
lzVJDlE2E5n04TSLhR7IJrkIhB1M/OLSfe/ek7wqSO2NGxIhP6NkWOLIulncnxfVFNxPo1vdhoBz
qgmAElXPwRL2fgjyG+HiayFTtRh3XLiq8/gtRkyejEagvrPe08V2uuz//rhnaap1Fsetae++VcIn
mR/ydRx5ZZKUC1Z51TCwqGdQsIEL9KspBG12XN+17+Je3ouOqT1OOpAEPqTmc4smTaRjo4NMrX9J
v+iFsOFiLuenfRvWUSDfioO3IV7W5M5pKykF8+GSL5JPU6naXxmTypBfBJZCZpRN355QVL8kPe2g
h/ZqKig1UYMVa92vGaGGtQP+TsvAKa+V1xUxtjGgnYohk1UfJdEphMx05n3ZDGU6RVIA+dyybwcH
Vz3HI2fZ2ziCNDTzgHqQ+cUbr/tFx7mZeGYN9ON8L/deznVF/GapAuRUUYb55huojx/CJKhbLUwK
/xpcT+p+aEFKbxPmNoaMDZTEU8P9dGo0qc5jSfew49V9X1caCRD8zCJSVdDI6yuPEjDP++DG7nNN
d0NaM3B5N0Ou1jTXDTM5IRAr/pAtRvoWwNmOhsYUiip5SrMp4u3ohjylVNp/lidBtOGqCkdoO5Mw
oXO6GBYQ4uKefqzsz7PE7/6v3svwVIrWzDeVTJUbCfPUs28C3ucUequGwoMgSMNbqXbZ/jQ1BpUl
CE1qSC7seNe/4Xn56A7rU1wLkxq9AdAP2Eq/0LOpYo0uCA7RpkcunEko+12nzxIB4kFybfpZIUAl
sk1baUUUtxN7I94dgNsCR6icJbCgNfzI1IGhMAAXM4mLMZrKn7YBw9+wEx95wz4N2yMqNlBJBsxj
ASDGI5HpdFp26mhXcYoM2OU5DG+vj+4uyakRTKaixGyJSvwc2Jsps2WhU1En/yX3n6b3oZWDSFJR
9JjDbBUq3oqWuJKwkWi06648MGzrtiHmhccTiWLFdC/YD27Wa1x7lxnqHs+FWKCgei59OoI39V+F
B20pXcc7Jok42cLJjWBybRFXojhZPAtLL+LuFggLqk/7s/V9a6eDams+xAiglmQrOyF9syV7uneA
OC1pNe4FnaACNRZ0995sWM2YM0/gt79VYil0o0C0OJkAxsNsd87aonP8jgHodaDVqCiPDnYW3GSt
f1XbvCMbNlEstyd/Ik6tmEZzwqPxwHASGWqrGSPImHxg2ic3P0eG9Qw5bETSxZqLa96mq9EXUMDr
wyogouwX4y+axzx8C7tZjpxeeOi4/eN6Xk9BiymzIABdRpMz1SUCzOltqy0KaGY9gnLVZ/o94Yn5
AXyTfPKfP+wIMHR4xBwOxLqFIEm91FlXTJs1BUxOLCgl8wu9xrFozm8G6j05ego6oAQxwFMdQQ/z
jhGzwDY0aXrCfzTlat+6d4lXKD6MwLdcCDAozHfEo08vOjgRw+oQBOj2ygFXLcBHNXvVYfz4v+uX
IaeR9CqM2arAvn60XIERHfs1OIPwrlyZUh7hYlb35F3i4yE7NQL+jwgpoBiSw/bEhsa8y7kPChWZ
rKhKSkGQlYUy79C08dxmJpfkxTvPo5s2j1YyTtt/wf4ZsATprEEZHloCcYeHGfe2CiSWHamLHGPC
hYqzvaVeUE44AcvrL/B5cYmAbFMpWPkbxkMXvLnHl0kJFWc0+HP85ZDuqx5gtWpEhVPoNg/+o9uk
p27Cf/LQwieC2ElA8O/LxF0/aARFYEv3pDQglCE7Re0EbB7tI1bS9aF9wMNnsMGPnTIOp8gURZKW
nFlNeq5pqo9/a95tsWAavPq1jEoYGMEPY5uKHdDWOGD69absHrSv6K94taNOduF1DnMRepetcEMC
4zXvV4tSMcHMsqqAjsjBzCdNb+lpEwIBYl/YLvjnytiYjTzK+ZTvVRdy2WeyWqkH4j8JKKqIB7C2
AezJPBZCeJPiwuAVkB8BEruXGIrWrWUKLf9LcyhLwD0eNEW57Oyrlez+www0Q9ARilQWQPeyN5yl
rszbbyKrVnn4sFf7c3iw+Gl1ufzTzPb4Dyw+98++2iRTaheF78JYQbHGSWs6NsdSS0vakl+4qOe8
Z0yhCo85irsoGl6mhfwA96VyfUUDZzG5zwfoscTBAW2g65TVSKlDuOzDKtiapamU2IPw7bjutT1B
iB8ZfTZmUjKODqkHzhdAkSGjBMhIsQU5Jcr8SSV3j41+CpH0LD159yzkqtD4orguxnI8DIR5mFHq
SLCvXJRvtolKAXrBgfXZ9t/jPZ+EovqaW2T5tpImtIlmY6slk5qRiZw9+uR+gEJvWYGNqmjpxxMj
ToYhvzge3qfomv9US6/b+1AgOG6Oyvi6sTMCnENmnoSw0a66hHYO4HvSyXQhSuT8+zFHX5WDTn6Z
Yp6fXTUQ1ID2gAfdq6O6Orl9MikfpdBAg91/vcXWdiBTuplVxTOYUuAiOxp1Pz0lxFIZGIUj2e1K
KDCWP0cTOv0ibr91dAH8MkANfX3hDMX6RaAeNvycusGKbnwFOUO0XypokicdomhlJez9w+/4K31s
LSPnTgt7rsVPpW4h6nX3ly66s6U9R7WxqMkLeklhGOgmA3If/wyoG4+uWNEd/a67GuSSXgM+zA63
y0ODaxvHQW+1FM9mdgDxsEkF28bl6mTFeEHu3fGYjozStQmvpXoAn5il+4V9sVnO3kUDtP0dNjox
nPnZCw5uf2IltpOsJRkc2qmQrnd3Dw0gvn6P/oboFMEFzZO5sW19zzFSu3PdI2OaE7iKhFWTW+0Z
vFat5gk91XYjemoPuaHteMPix4rj91xM+w9dHK4PkzrFPFpj62+frWYECFPlRLESlBT6nEr7jzTK
TXlgz2rW0Nxw/OZbBQzlDdNg/8yia9GXed2zP7HwMkHMb2k/zUZ59s/upxOYdk5gsVBZ9V8ZZqdb
XjM8fGzIpVy9DaOZQiQ1EbgdP1UPVJiYwpccL7OS85lgrg6VqW4Lv/nhnS12PQ2jFa6zZP0uZxPY
pnPF+jFdHNIPCr0IMN7RMNGDow+mcSHGK9r+KNRvOqkD6I+H/C4+AfqLKzWBuyTg75mxcxxwaTUj
BvQwfAI5i1KJZ5PuVup2R5iZgimrS53xj+mckoAJVUBPhR/jmRiGiETDIMn8h+LT15CiiHGlmL1t
BPRfZPDBZQLHaNychMwii9b1QvFP3DSlK0zIlme9pg7lqcOYFHd0YxU8/cookfWBJahYyiL8Pva7
iA3UwrHisbP999ZabRgGCe6O8z3wA47wglE8oVZQAL9oIg83j3U3umLW7ZqmagJgfy7BuUey/RMK
A2PecJQSUX6EX7FZAuVdYJtPBwQk/3JKfWu9FneOKNELqriyVC8riTpCG/hQ+YLu6oKONhTac4wj
oNYhPhf8xDpXZSAIr2W7/IIQYZY9FX5dM8masGsDUko4ClMQnYOEsKBeMPLJe3T+m52qJaj7ZqFV
2wefZUws5ulpsDpA5Sa1jwHwmKCRHcwkAfIMLLVeW5jmzEFvvEarW/eMiTMtUGch+a/cXZHdYcjW
ugX642tdOE8KMkMzdRLI/+pdBGYYUmeKSQjL98g+K7IhIE8t8xG+pKDvjI3D7s6EfPRdAdKcmRF7
1gRAf4q/jA73AGawQ+ZJJTzUD3PA0slZvB3IxNeYmWT1qBxKsL+DVSJCwZsL5YlGN+RBuRQwwVHG
7wVIwXwRMPf0359+uwskXOC3MKKODaSJzfybnLptLR9tb2iKJh1Zqdqp4v4eYeaef6Yw0E0H9QWb
wQzgYyV59nGU+VBkvMIxHpMqvW+Vmt9RfBTNXlPO0APXQ8nf3J7+1VAANeek1vvT/472QEOM2ePP
Gu3YpymVMYbFCbwoBWgGOhxwz7u4tRPekLhHGcYpKS7L9Yefs5UVGbnAnFUgzXcE150ggyezmzXU
Dvh/BEgTJEgWET9renN62XBZ9xDsEuTGaN9jO0OQdWXuj4WTi9s/g8dFMlePmdLs/ONY7js9or9r
aOUMYMiavJtZ/71WMNc0O1GNZh62r5ItSfQysVLx6qViPJAkZAM30dM33M3SVjoo8bp6BbtPc54z
boqqEGuyu46PInibtt+W8RqY6cv91duMJ0n9FZLMoC0XYQEkpyvPWuE6YT/TgQUmVfTyWajnqC1q
3txgJzfivdzYa2HfU+qoWk2Rk+KEXVX59GlA+gTKVqkwqVD393H5yWlQPsFZKz/GOYbpXzbGlOPR
QZHGRRPQcF+TAm69FaUDJAVO2sJigr0YT6GUEx7s5yXK86EVnDhUgeGFgxmPNzEXVMrmJKkWtti+
TkQFGuv9BgAGykRaIDStPYZOoGRnIGJLlLVpM6ECk0/NFdrBcRqK7ZPKL2x/6NJ5q4BOKV2wEH0m
Bkw7t1JR8MuLkbk8UJ4SmXA+5Oa9IeuhduihmltBUn1yELKvh+o8ErVKEqAVYbDGbMQp9p4aAmNt
NIR0vCUiiHzsVClY3WMI09WYPZ2rZE2tASUXSh9LPDZ39fpkgpCkuoRnAZVGTvLvTcH2HGqjlRb7
eQ1MfVQ660m7oQ80Ha/lYxWLam7qLHmx306r06p1pJNAku3qd3/uHv0KNKlkCx5ktlD9aKBTgUsC
VNsSAJwKP1Qo7aVR89US4x3O4pml0HbjYHFA0qWEnuKsJ4eoKJfH7ocGYwgIlPzRbdNtEmCCDHXL
FhrqR8Ze5TGMx9Bf8RBS6Pm4p3NZMVcF2NQM05bteia6qFdFrQ6XGTXw5AInAcgWOlCLwjm9WNrA
IhTWUnW7Y6orTzGG/J2Sp4YER5oCQW4vTO/HjhlLQC27JfY72karSj4KR3kPPa5ykUGaz2W/8M2Z
d/+j6pseNhJAkdkULimaMOttyO+qtXntazCHcEsu8d9LXmkDwzgGaCFY5Ib9Gn+2xgaAFIA8e/m7
XCH4/1LcYMJtbAAuM1popeKXE82/16jCKLXxiKPxCn59EZxXdP3mlPrY1TyLG8+xznCOzxSe3WiE
aHoXmuB4NIfMviVntsJLWdtN5+xekf8+F4Xf37FM93QbUzs7LWME40JG8PIaKeHm5dAXk8pffP9f
bzTmuTq25N8W7dxmSr5tyhIZBNqt6kaxbh3lM7ukA7zDCZP1C4YxnUJ1PnRNwllHYB/Fda1U8tcK
ahSCisc9Kz8LpqS/C4DqgGwEPPygvG8R/YPIyc/iVTqjqYpKiL/0da2giIH9myrmttxbfqO6lik7
8RSmm9IsmNgCFLWAkJSM4clTCxVpyXDChQdNjDkivRxs2wpgW4UksQ17Yru1EhqTG7HGR+AzOAeb
5ThcA4d1BQUXgbtD+MFdmmwoJ4hHu6KRUcCZAIbnDGkdEHFvQujJgSsrApve4iP1Ugrek+EQA5Vr
8CFoYng7zJB8btYHG/G3qYaVjbj56BHwSPGvjfXseUxi0cwzTPafPv/6wtUFPfeQpcDhaj2D/fc6
Yw8ktNzNpSBmTB0ytMXA4/YGzz1O9SE6WtkOZtA7uGS0zOPlwaNOKdNE2FCbY98+xZ0VwsjHII2j
tPg8jnxxM79nnUy+VGoyHon5mTlGD0u7qo2a4pVlfJhJtRcTbDOKOkOJrNJ0xgQY7zS7fsqGIw8u
eiA2ZtpS6EUu7Zcx0T2eQclSSBOrMIWAY4nNCp5EJlFdkJ1zFgQvX81mWQdUPR3Mphty2itg1nLO
RgttDr8cZOeScVKRWPrulamuTG0MC6orhx/pzbL32bGyVFO9HXe3HfgBaFOfd+NiC4raRbzWfZAa
fLvyr4j+7aQ6aqDlb1DLjOOB2CbO+hWBy6uegYzRbJ4vbeAGab2E7d7jSmRfO60GR/xCfukVgISG
GnnKv9lJW2Z59/oe2532IoKTG1wNI1DMBxHZiIjb93CeXYwb1UBWxSO/aa5g8csjq4rWv1Xw6czs
AO3+hSzAojDOSeJ6zsBRzi3+Bb6zlJ1O1aG1Os9ADkBDZv3FPJlfo4sWfdbUMa2KaJMECJu+eSVK
fwrOqFfr4++UsJSPga8alt8k1nCQEjYieL7HI0cbBE9lqSpMS7CuBbo0GC59NcXu1AYWPbrj2Sxe
ykssj1hsAOo9X1D1hucZsLFMG8LqcAI0DsQACIAsFshR5Cn6R7f1B/fYq7JfhC58gx3QPSXKTWwH
/noXLwogUg6sFAp/6ggif9ZSInJnELCLnRThJ8q665QPe/mNpVItzyYwHzy8s6X8uQn4dUIK4/i+
ClMwIYqDq4NdpoczoWIjEgAHhiqjUDidFIhbEMF3omJdKmFz1LlrBbyCd3ff3BsGDvMWP6TQmt1e
v6e7CSxFuSdUaw/kqZN5PRxDho20q7JY1BSTOI7vV9MCE7WRrtUlMK041dFMwJMeVQFuWCogFWhA
beczV2cfH9MQ7uhxL8Q1gSNokY/tI+0vM8MGbHKxlgf1FkYUCq2SbYwG4v6nLrJPwu2ccM2AA5/F
FkJxCGsBX11Qs38sqlYuN9L3lw2mSqJTKOcYdkRYfidud1yOhvuTVp37xL0M17rL1CHuZogaj9qO
oO4jL9l7IiOnOiCrv7V0qjs1co+dKy1soVzyZHOGVe03azTFD27BCuOyup26MpyDG4cr2V5LrYxi
Op24mP+6bbX4Yz8dXrnqMM/7e7pUDrcc+EpcBsFFhMVOF/8gQZ+dT0jHXRppmcse1NUqvJ5iVJ1z
rpmi1sM2uhyzcXMT5Eozgj8Infgxs3gl7loHB4Z7UcuTgXNpNZvO8NTzbpPlhYTSobx1a9UvZNbn
WoBxdZUjy5ocIL8/xZuQobBC1bybVZaVTGUOoe8K6JHIlKwyq+E4jkqtsok=
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
ga7z3iGMhGhga7TzPGleypVOHJn9S7KEP16RJ6j/y4QGRddc7/SJdXJ2zPvm8FTCqWlJhu6/s34X
gPP3kw7dN1YdiZ3wZ0Vzt8uhC/B62KTkMGylsJT3Hm/4AVsby+VuOus10FHgOgp78G6FqJDW2hD4
FEF7AvpJ8kF9S1ZR/yBaB9R5/vEzgMTG6H0b1hzTpBGPyaW1S33KG60mDs4uY1wSc9WkIOuDsX13
gE5v3E3AdV0s35W8mk90srPFan8A4v9WhQvKv0pRdTPwajKYNoHYw9l0a0ijfdCCo0SwbSJr+KOr
7KJQNnQdeGn2Y8dg3BGFPO1H0k02bZuSqUQ8rQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
dBwrqXpaPIvc4b2fzIcAYNKycDBKm/hw0N9OirP+O5J0w47WHpIJLrz+YZdtlXZ+W2OT1CCdKga8
l9q6LpHNXfMJe0tSBaUQJS9kx12QCBYd7pz6Zz4XteULmwejqAW/r/1SNtjKdsFfgoOhPbvsYv0n
RR9WE79+rnvNSo03sWloLz3If8EsTQUj+4AuHA6W5eeLCFFrjEJDELred9ftNf+GjbKQ4DD9VT1l
GYpqKI157tMW7VzaYctB1tIYsZm6N1scQY5/pen6aJE9XG/GVJc/lUhiKfjKkAB4R0V1b6xO6o/L
Z0CvpttfY2ekIVc0VuCKq5gMTfn8BkW7RjZNRA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=9072)
`pragma protect data_block
K9c9n0r8UqSRPYbCShNJbKUo8nMlqX/ARUm1/PxkQhf8vpP+dVWxtXojBpVqC3lc2IJNXRVs6uXM
vneWn1lOqZ1DGaGsexVzKsl83EBhS5FXuFX4DMldc4XxE3q+spN8waCJ2Dw8YlcOz/Sjd6mzHUvY
qZJFkU9+AIbmwUxrCrlgkV/c0byGARFHwCFBXjsquFfamhzS73bcV5YK8GctPH37nEJCr6qgRqXH
TzuvKyx0JMExZSbt18XcEBEY14Bd9wu/ket6kkWHemRty2jaqAjTMaOMr2RgJOfIOdp1hSTc7nEn
t7eLEmCeMvd1dLvcQpWDIe1LjhsicdBZ+hXVrZlTxTeU6Kw5melaLjfZ+PfviS8Sc/aIRiXeeO8U
5jqojK/I+rwpHKKChUjPkJ8YstLhQhgEwpxhWP4lBAt0zaC3kh4R4Is893xLW/mFPoKowKoYRav/
gqC8r3rssAGSyvtURmwvl72p9y3nH7OU69VdHpxt6IHdcfB7maVpXbcZpSpNU++f8M+AZO/fQ6Nc
jap8GG7gbPBcqEogecLbmTVEfmQ5cj1R4lcDOxLE82/FgyF9/TkmE4/AUtnNdvE+SdiocVdut4fT
U+JL3OLWpv7d6a9nBS2ESODnMqcmEWrag539RwZGtCvQoGoD7jfdqLESZ0boOGknjA/xIvOxVTXW
CMSbE6nKqGXu5oRSk805mGcpMOJzcC0qUf33Xh3OOEWYPHoqCEANWdZfWy22mHXzuobGuP+KjOz5
Jrg93M/7OUOlZ+9zPqP1wEB+bC7gHoEygl3EpdeC0m2fXf4tz42cadApidPwN/FVzIoDaFCvz9dZ
0k4mEAjPyC8Kb+7c5WtCqteuBeYV8AsffXpI1fHhMkfw7eM+Oo5LQK6ZG7pzl3mvjTx2KfQecTl9
w8e03kV5uNkcd9z8b8p3UXq5eVHUN2C4FuKPUPeYh0iIN9dLzafgfslwEqgXmvxItHw9yqeTpaIf
SOnqGAvpT6dcRls4o70mGFrAZdnFcsh3wWO0e7mL7QbO7wVuT1Qu7G95Gf9ZoAQuC7EqbZj5IDEI
0SpV/THnlHTKJoAHrTC2WB3xRcU+3+6P6e9NOgLj6Lm3CaSw6YKLNVU4z5Ydaiontpc3+UXxey5x
jm1oYpjdGAAEoZeHpTgwC1cNYzq5mKorZlRTj7aBu7RjaV4dE3WhT9JZa4jILY/nz1UYk5SroJ0i
mLPoWCB1IzDnOQHbEYBrXS1tJmru3vqPik9wOGgytPWHnopUYbIDAL8CgAl7K1hOAcbNdjr1wZjA
rx8XjLfzgbEYH6OoQ+l9Xhe4IlgJZv/Azx0omj3IMjbjcZwL5U2YgRiI1s3W5UCsIs3qF4/9LnsA
V9C7t099xVWYvS44QIjM16T126nWd69g16zyHtkA8Sl834EPxB3Pj52TNzVHH0bmC2CmpmfnUWCb
4Bq0kGdhLFZHfR2/OWsyRCcf8SGp8bpcjduOHiGKZyqV0xGzhw5OtiRPtqnEnE0FTELRDCNyWq8n
s2rQvusBd/ClRE6RieBXLASIHPo2kJWBtGaz6BV+qNT0RCXXbZuFKrNIFbEhwMOC7W/BaZsA6gxA
2N0h9GNZvFPqdrbwHWAXtwQSZ0puDDfSu1M9XG1uNjrC1aN6lIHUGIIZ2aLnsNVYyejKuczoRCBt
fpRxuuZj1pk71Im6az2Vq5hGtaECuUkFi7PhUup/FqlElAxVOhz/38wTBk8d7yv2XYxi4PSY2WOw
ivra/S0ZXBw5zdiy1cyrw6yUM6Y0HjKXqHNzRkpC6Eyl5z+uPneWCDHDV5aB2w/xXnV36q40KopO
lrQX9KPda9MDau6/Au2vz3JHrnXXnJzuAvXSsWpYxgrfmyKUSi2GGL4mHpY4bmARGPo90i8YH6fs
3y0um88mF0z7/HjxR6fmTIJyRho3QqiA0QABu8lLyWawLQaO3iGvUblbHCxXf7Pftdju44DchqGm
rNJfrZSmrcR3FDuJImQ9xdDYNyyraqj9C7eHwI4Pnems7Tu/DXbPdMELYfIQAxH0BXNUCV492Ala
viBDEGTNoTkS+Xwuera63sI02NOdx2nkBn9shmx3tDJuCOmo/Rr+WrzhyHjz600MStkaIZ6mW15A
k2eCUdiOxllUmW17BWrtwM2FAtLFl4ApJELjb6z70GiVUDv7ImRWzdhyLiDK89H8D4/ruVCT5+AN
Mtsb6EshZxUXmgvSwIyRyxfLE0rXh5eTQb4148SO+ABOVuIxoo78tjpdf/OlyIuUDUIubDgJA61+
umgZ7cluVkR4R952jimHUa7TsS7C1PVst8+CCBFqc8NLOyKJOvv0PkRtWH222Ma76EyOKqUihOAP
cKCtRDDHr9kiaSMl+hHT6+ighidT7tJGypGHYQQkecx4ioIFYOs2fT0f8WyIkyhKt0TEPxl3x6XC
m+KMDHxEWxrFJytafpX+j2xsEExe0kEJaNePoAv1uCqIKYCgBsoVaBZahv8zSgopqmW5iAjOnSMI
2xu0RoM5sCnORR14x7ezpIKrUV/93hMQgREiUF0kWEktwCQJCwX5ebtYP3SLxEaW3H7AV9tnDSe0
De2IIxGMoICs1rNwLrig0rwxPh1+/dNT1h4iNbssEcVQKWSM5Xuz6bU7C6bba3pX1C/WYaSLzjPz
aAcvSdYD3Aebaigp1u8vGmHF8kk8bcjtxIpAOlBpJhi0wW5JhSdbWl1q2AGitQMxY9m1n+czmelK
d2NwL23zp4DtGb//3eH3aOM089WyuPOJlB1BJXkqzClxdgw0LpOzN8uWZlLV4XGgMDD6XdF8xAYT
zGByvVujcf3MuFKAIR17f9oy+hJiIizJJ+A2dp2ewBkTu72/aZp0aZb7ZYHNOXdxfmgtLXQZRkGr
Rwu9xZfyuR2RzcSBHufvTMn1skonjESonms7CvqxTiUxRrxdLsM5daqaOr3nNjoL1asWR4nAczv4
zpNDDjyoGMBAUSex3t12sOXUJaTx08qRaXAGZ9S7hJuopUdC6vWP4MTMZzjlRYxEy9LTvcRn/xAP
xJU3kMsY1CSdDbZj5uH7JDIls7WZVltAVKrMlwaPB8oLQQWO1vr/DOfhOTT2SCo0xd7xVthjsxFv
aT3sz9hREKaNtywvW+y09vdnlYVRiYo3ONN8yOboqQ+JPaw+y4apIUlW2siH+k2BS0YXKKe+rcwc
R8HM+Azq8s9svgxiraPRvgGnEckR8NBkWX5uGN34dvvkLoLvc1ILFOyQ/51j9H52rgrHLZd3SUTN
BsYglX8vQG8AiQCJuozY07ijrdTOyyMX10NDhRFc9474Nj3/7uvpuR1buMO/Fn6o1W+HFg/Bg9C8
01j6nlyGJcfbjaC2HS37SfuyjoOoZckxmltM2/omN3yk8JSFc2O/mBxew6Qh+Ly9jfhI578MFi1j
nx0+tRopaWH7lzFX/lTCcGkr0c4z33HZHbI6wjAqg1ZJMv4qjn9BWwQyK+8x0wJc/UGFjrifDfNl
9h5/UPp/gXAYovAWHYx+rUsFrMgyBm6oR41gppxue07IYvDa1ScZTDE0kaqYXCWErIe1YbeWhEQB
5WlcLwsQBxl3P+qw0vyU8aaYSdEkTSSQFxhVf3fnRIkdLs+M3juPnEGqEno52882OUf6K+alt7OK
Z1g5HuDmdOnTMMY8j8PNyWU/gM2x2IMxNSYZE9464FJoX87p7KxRT9pQE5A/+EwtXRTG85YYTg9X
cNddGpph1x16DuHqMYK93rjWLPKBQbhl0XkvKbVyDaSdbVm5ZYMrUQl8mEX3803f8fCY1/HPJfQ8
y08Tk6tM7fTSWw+EM/3FFsqc4aEBU+++znUMd3BaxXgEJvsxK1wTOJXlMmb7CWCv3nVE1cmooOYo
gUW+tg8RHOTVIrNsWRpI98hU08T42UPcYsdBe3XFIrY70sIH1uoOgAmvWihMaVlI4npz+VtFNwzF
jbDKJW3m5Fpu7uqj7gHc/LLOkxBN8VTPscAZ0JFqoPMtLLZElVx9/gHWGFl+ZtSpVSk5aQ7HexxL
PAg0nfeJ3s0nvFI0mGcai+brUI5+P0ByuGyu93gDpcmz6gMncv+y72ouXoTbkoss6+GTJBkRusiP
M9tgwenoaO25M+CjCER2B8FkfFjZdij3vXPHrjHiyKT28gjoSJ4jk7x3ysh9V0L8f0zP1AFS6jeX
68idF3H0iVduzr/xdfo3PfwXnrAGOHFD1f10B3VZZwIBNBgkb7fpnRnzRckwpTV3F62QP6mRz60x
wXG6t0S/rPhBtrAtmHQM0/YbLnkJvvdB9eV1NGpGU2zm7lo8+NM/xXsj078q6J+c+n1fg0Rga58n
YWVkCrUyJsauKFA2KDo6AJ+f479Rtit+fyjIFmJYTvbtUlDpZpdRW+IJ3d5b4y+hCt7+9l1O/+j/
jzZzHcQ343zUmWlF0F2W9onHgeQ6RQ1MaP7kjYdbyLFFmbKYJJ9cNNGeZXBhna0eZErEvI2XaoRu
xo3xuDVt9MmUIR1LgqndyTWyOi+bWNbMekvQf2CzrIxCU/QOhd3ImkM5RrMrLte1yVQLTZxzNd4M
nnsuVpi0ESJRQhkHzssP8gbNAveLrV1Vs4o1KIF42O7TB4SeUMdLfLVUGPd9Uum7rbgK64KRRi3t
+G9iA3Tiy9kFzX1MZP1PijTvNUvOUTrktGNJ8yIm7DG61H1QN6lJm7ynk13jzUR9nRfiYfOXM9G4
ewXLHxixXz4/54orK8TZBWBW7XVg7IfZ5QrY0m+elImbAzLc/Xnm1OpxTh7kgS/vNptwwbk5QH5h
d/JDREK2X9dNZ9bAqA+jcNrcyml/oxOCBJSRctWrZUciAPJzLEgGSMYX2pgaO/TUnkMfrX9jM9Oq
52AOUzYJ+irgidgbra7jeprfcSAJfRekv369W5TZktDpqa+JHX+D4xq/J/Cs1eOiE0O3QzhToJGx
RHty7ZF1BkmN5GgQjN29NZlUuWPCtdPgUcx/j7LOG3QbCiVbNl1Swb/+/CWeehtEG0KKic6RrvWA
ecXWEMF+6WjkQds84jupYBBJbk3z5B1QwOdotCDc1S4GE4zBcsRV8m+IytQJpI5wYJQMqyzCVxpV
ik2UpfT/K7xfss1O0zbxU+50gZLudlfPAHu34vH5RsCwko3JwMxqtecQDyVKJqjcemc927oh2BFC
PWpyQhjWrNO6TkQnmIF7mxJiSBR+rJcMQ89USx7CO9g6dc3Ml+8RMqi8teLLDE41isKaxqR7QpJa
E75VlyeZ7oCnnR9MmI/AmcqZtTeELvW1utjYjUe/Uf4QZo/bdur8TDWdrndCGMcBpXaIjeEIYskq
odTpTNr88KNA4umQ0l3SvAN45vyZoOYkfifMF5cYlX/A9l4SC3MYGkE4cdtPB3fzLAiyDjds3Nz2
RsFiCBMyuh9uy1pcDZvGWUsB2k14gKKQrjsDw6OrtnAaBD8DZGmEh6E5yBPv6wF4hX21wH0pFfQW
/EwyNPz8t1TE9IczAmyBKuFKj7Wlv0z+xYjU68C2RchF8uOUsGJ85l8Drudgim0V45zmdfRnlF/s
xZPti/03loTy1iDH2XlEwAQeVTKGJMMp8FR805Mm5+CzbS9vm7rT0t7xhpJ+MeR+4fSQBS0e98fB
DfK8fpESNNp6AJCoiuCw8Qe89Ew5IqC0QN31ABocnkyD2pq7BWHs+cv+tAUk74prDCYRPMdga4H/
hf+ywNk9TTAkqAGSCelHDt8UPXCHBZ1n6dGuT4BXs5EKGbleNs5/uG8asjzjNizHmSqTqSd9Z2UP
6pDCeImY4ltJtMQGGfO+BfOJcd9f2B+ti/94ymvWf8z/tFA47CD7xeb7EfV4w1gIe1Tq0HWrCfWh
s7ANQHGFU6lmkdhwFTcmXWQZfk+yoeIBC9HbQvcCi26Oj4i4zSCgdCbJ3c+OOJa73DS2SaKJPewx
hGnCqCHNerldzey9vkTRv06+kByvcMibGewfKO0FJIvycqeZlU9cX74sqb/ShTzaifemmEpqSGa8
8IaIrwRATydXr0+SzV5wG/jeJaxVSf85r/sgyZ5KWYNOx2IZI67X5BU1DNJNYsHhOXnL3tFN7RIb
8sf/trb5M2Cpt+9zGc931VDiK6OzleASV9JcnPXpfLhya/tzeYwpimA7PB3/6BGbpQv9LSKPGe+R
qKskLMJf2Z1XBzx4ZX2uOAawVthpFUkG/jyICFyKRNI2og5V7EyaZjtN46rgvHbIu9Fmlt99HPpK
1RWQvIFWxY3Xb+hMKumDbnxN93nr9pERpepXWoUM+aJ5UEfW1ClzX0bDnHdjPJhlzzMPVwMsgisn
JXzIeVkqfdSsx/6WYvKboo/ozUkKDtL5AVDE+jeuJIg3zfdf3Jkz3SbHdjnRoMIpr6WoPi/ZHza1
uL/KB91LVbHd9vXWxh5HYMryhtQxhg1QK9BRLiyuzzFj9sa1tPj2fcv6UbdxepzuN2n63RGLaqpv
KWNQZnTZW9zTDDqAuirGyK+y2FehRoutsomg+CPTVUMZIp7eQOCEc260idDoJEKoSzNx4fWwD+Uk
1eSTzMVVdD7lImjUz0xHylKL5uVfNExQST+XZsnCSYM9sWhL74wsxwg5I9gJ/bD/NnfeYkUpjVpw
gvFtr/fDJdLNrbN9sR+tHmyf3u6gnV2eukNw3ZYSRmrYAR/7D3XuMOG991WhivOJ8h9MTK0uJ/xY
7u++UW4tC77/8Lg5HHpRUM12NWQwjJ4k008HjaAaEUHoJkTyNYJPcCDiBv849Ex9rwcezlLlOV6t
GhD2ZkpZ5tBo6/T3qpswHlq0aQAK8Jaup+EN7GhIf2oNJB0jrYQHOTUoi+Z3PDWmSyOmnUHU3ljS
QbsMGXicuGqcgcviCzB+xK4jgMV9sSfiTdeZ2zY2jlxCYTQV6y6WrjMJz738VWejEIX7RiSWx9B1
mXyQU4YuitlWUGdP/gEAicJxkA7Jp9lKCazDkazXoC1qiHt+NUZivlgC77W9wZPv/cke4b8yxEX5
lDfis+B4w13hx09ffILJonK+uVfshRxs4bFg2AuilbyapdI4+rcfEjSD63b/d+92uSUOnDXIZtnL
ROND7DR0be1cvmVuHoBrC+7Aj3LbloDirZuAuXlNAtHdag+y/CqeLtDB0D+cQXI1HUxEvZD2MToC
NgHnH3IbjchGQzX8VAX90WRqJc93/X4eV9kgaif3cwWagm9lShW8BUKnVNmb2RLwq/wk5Rt8kdfo
Pxac0muHdo1egINWqHLSlUXdFHPh6skoPuoAN51NwQXTSj1v0uUS4cTgGsf/bFtXK+SSsDFWc88y
V5/twDHKhlpuf3QfExNOWSKtOHPvxi9WZeA8wSy23wv9SPuFxKaGE60AL4xn/n14KwmPSn+QOxt6
Wu1dAsNbYut4xf8fzBJ7oJcpSYXfrk7XeqfuAK7jgrA1piJ8T0cdCiUuveViS1rsY0x5LortdEyg
RIG4wtgTRGlvi9lVG3hYKP/2piLhQ9LUir3lG84KU5ufHQcownlSahXPzFdKiNqG2LyhHJjXnQ8d
eEE2OHZ7cOvvIparmWgwL0MHc9Tr90foa1+MHyOEeHzDPytUGMDSYMW65ZE1nSLnpqUX4g1BXpeq
oHiM83+brmznOr7C8iSeAJC2LktB2jGaDNmdNhCgYU4t8xNAUkHZ9pjs7Hnlo/Q6UeUZSE+UoR8w
Po8PuS9SAJI9cvay/1F2F9vqnxc24GiOhLZy/PROy7TFpSBG//0h9nP+Yb2AmFVWp0+UlFaKIR/9
oZiVhPmjXoVnh27P8b9lXxvzoMRll313/Q3iVYsyjyCZPhJrRFb3HKN/70tlr6ZkLlM8DZVKmkTu
MGN4tWj7cKxFddtRzedRRo54DnxfuT2ECIWFWtv6miBma2/VBDTtEP6j/NDarTtSnezV2cgETkmC
Wk32LNi/5cAk5W+8yi0N5dpNInYYnD8zuq7mzfWw9Pm9ViCtldua1N21zNUOW5bxfZR3p8P2NIBz
TComnF/9l15l6wKRFGvQhh7nkaGVc2LQ1jbr7Mz+PCKPhIggLrzfg69+rNA99R29zEALdx/VURWk
mR+56TPp7tQbDZLpnsKjolicIVk8S+x1xIUnxFdin6bYDMkBXjqYGPcKtl3niSe6CMhFwWC1C0fI
S4rkQq0TdwMYn9TQ6VoQN/WuEV5kJDDRBLFZBawUqEyi0nLXbmHfbgrmXlKF2k+3k2Gfx6g4sH1s
9jIdIGZB56AAQSQEb6tky1HlAYK7m4+P+XKFZ6PdRMffcpGArc7SwwqErQGNuUyQSeF5PX0mT+NH
3ufPvO6az+Ovt1InYQHtKKlXYBt4mYSB9C4e98th2gPKIDtXPVyKFzl7yIEWAlgyQvmvfLVTUHww
gNMo6qyH4dEK+jaI2sdVXWrjtTkfk+mc+nGT31Vuq5tuVfPq+cBnUPW6EWrComfM6JZTfOK8OXTP
lqEVNbVlQchPSxf/8NKWwzmq39ucsadjpJQZ3SwBL5bV69oZn6WjaR+JbUr7ui6ERBlgukdLRbOy
TYYs6kXOzElrZFjznvjwtJ5dttrKICV3K0zSVerEw0lo9Q9J857OIAOa+SN1yHTwwVIOzIlI5ENO
qbg+G0QyFuMa8QYkAwKvgxIcy5/adm2BzUQ6zJH+Sd3+l/yARt69TBD2YjMmMOAMNJe/NcrMdpep
hgL9tMHzGt8PLWlfkbotPg9iUWtymbpwJ6f5nRxcVfWsICbc5OzqDll31ZLtCPYrnC4MeFsbBKj0
pHJouVEncvBLAKDtn4yui3QpCSKQEZlbqrHLUmbnBqZKeBET8puoZnDCovKxQWYaIMxA1F19cDI9
j9ko4lttHDGADIgLNjApkanfbT0eEM9AWFY4C2IsJQJYoD01VhSPuQyCnshw8VpwCqHZyTDEe9fc
il2cMe1Y0sxpD+mam3T+UG61A/DY0xv9lwc/TzeaNZByytk/J85cHBmsA98xdAih4rcFUpLkvpE7
cpBhdMuDs10EK+MDcTgK7ETwXDtVVshqjLw8swKVBFUyKteDF4+TRwJTvcTs0usj4CUAwIbIr+90
0sJholbcCFB9noJyDfKTIRYyHlNrUtc3gzTYNj1+GU8sy27CU4dl7Qdmh9uYTTh+9FfMh2jFzKJW
cqjZ0vK+H+vwVfNR96b7JXnoxF0tYn+3mW3qWtCpcLlFhP9GUyhHNaGM7Gqiqn1I1qY1STszvJ2Z
K5qmM+4eEUiaW7OZ0lHSiGva5+ZvRd2JCUTho5a+0WaZMT1OwSO5g0f6eSDiE0Ueta4truP3yvqn
PDm3aI7czjBGPujf1YGF9vrO+tB8Iw+wnp36ToyxfASS3Hc0kEl5nHYnPId6tC2E4uFazMn02Rzs
6BMtB3h498wmoN3ZV477ptA6CfX0oBCFNLU/9rnfTp4w8UFHIHPEx7P0LK/ML4gYO7taq12IDowG
e9N1EU+finT89B8Z41ORLaIVbqOQiis4mzsp4YjOkUgLRa4FRkcOC3tx76Qj3du0So0WyUZgFg6d
Zr9k8SkKhgziPGTY9yG/QlWooiO72MXeZI4SCzUMi+ZNnxlAkdBKCbp/Jwuq9AaR/snjuze9p6FG
e2osy4XMtLYrpjHgtw/a89vTtxITleXR9+j4Ea7Q/kbj4Nhqo818nZL27fI3CUk1pIB4VucE/bzX
FysazuP0toTXpTtupc6nwAKazwzDwigfwv4p9d3ljyndOSHLZDJxQmGd6DG4HpjjFqp3PDfd3DQ+
1xbGIGlZxwQ7nKyX2lDnYl8Brx92hYtUDFGV88OYs3eyHT4+1yFp+ucYhwQlTwrGjdlS+bZyOJkC
zDRLbvJGt27D8RjR5TVuJn8IrHwxbafrIHRfd0ciWYoxF3auLXYwLutKGoMXclP0CMRVHQW7AyZG
f9S/nYKYsheYU+Ij+Mwhxcsq/UPdw+puVd+0vILbnBrJQT4aGZXf+7MHVPlL0XMKBlaoBixpePyU
akaZgPC0AaiBmbyzdzkV85QkQu7nE/Tj5c+mleXPc7f/aafvszdjvc/lfWsKiYwgYo22Zv3SkHz7
fGV3YfLQJiTwqjPHZqiD+Jqmda0fmmzXh1DPYoI4uCAW3nwHkWIgiw4/1voVTQh/bwEFpPbmmEwU
+GkrGOmLt6HXUvr2UfnDgzFnDjSr7uJXXN61WKw+ez0XJzRp8QU8t9A4H3kirn6KXYw+IMmkNIO0
o5ya6A7IDASKpbKGShim4G0VRSc9IW/pu+s1u9WnynfIn2M4ifUrcCU4A5NtJdy6JMMS/NNVcsA9
h6AlNKhBl5On89zV2zcDP6L22lWSvaVUGL4DGx8OvBe+VCLoibpkwgQ1o4s9CqaItA7JMmKSxQNm
NwoN626t7zn69TtEVU9GpZxbow5mmGMiFX9oBL8YkJXV+JRKR1DYRpdjtno+CTwfi7YKINrcSnkA
VhlXjjfWlbYolHqwK7segvOQXPQ3hXu+Wsezomrjvralhn5esvRyBIdM8gxg2z/f3QRebP5PKOc9
lhFZcDTOsuKJTW7RjsSCFLRaqzbYPK0ByYX39Bn1DXwDgIZHWZIHfuJHNBYbQAYvkzLviNjqAL7h
tlJqy4qDw0HqzatqNTMfv8CGjiUatlA866OLtpF2jEjetLzUnEqPiGCVoi2SsiaK6tQaUwmCbpjb
FgolkGd2QhUzAcGl2DBeamw+0QIJYXHCmd2N+6cHk7IBqEC4IWgaH+erMCsqt9NEOEazzeboIsZD
CxykhO3GpzxS7p62dy0s2wlV8jiOaCco8/LUCZtBWFmK2X2qOZ6eWX4JQS6c2C75d9LU9OHRvU7h
GG/nLglBKuEBQVcDKNtg5wO9MH+4Qfmhj+nVNpbJfVr8U9x29hRj9Fi15RLMJFX7jnX007eLaHyG
a5zYw8QFW56Pgz6D2pqLzgoBvtT2oNHcnasqCDalXLUnOzx88Nk217g6ey53NcVNftv4mWV9YV5t
7k1/TeCv3Z62uSGizdV2jqMCAHi9vyhEwASxEn7J4NwewZrR2M54CFyfSXQbWIOxkItW/uNpX1r4
32gSUuSeqjZrqPaljPju3DX044Kr702Gjb1XrShWQftKMpzc26/p1ZpxQO1i7Vy0bsO+jr5VsAju
b/wnm2kePpfSR9rzo1rIHmPI34lrUJWzNEsIpQKWpGYGayvBPDgZaA+WC8xAuvdAMXgvFRlPG8f9
xn91ydEBIlobHteN6IeEaf/zgidUDUEBt5KmyB6v3vefRMNbVpOpvsmZzmGXPcT9gIvEt2MK3Jr1
wSVKsWRa8Zye3bE1yLM4OlQz2FbxRSqArUfUy9CrqcYWKtIfV2sgqrPohFV4HjkzAxN/4waLpBiK
Za9jKdK17xOU7rI0JsV+QxPN4c6gxohZmJLkhl7hxw017/t6S5a0gO6yamlZGJ+pC4tKW93I5buw
1XKl2AMQl+8nkGsg3VdxMjPR4PGfRUpgZp9LnLaIN67eePJuediBbHXlWcC8IcbMyCP+hpvsRqAv
f6XoYFKQrc5sL5HZJlsGQ5S28Do4ybQBgen+htxd/OyeNuTGxVK7T6+QvuYDL85lKigGDoVsQjEX
WkFD2X1KdRnXF9RicBEe4d+/mJJIewFMUu+ZK0I8J528qjPJ3CYVfSz0XsCQMI+176D7IKmLFA/N
42i9cEH5x76bSdcAmn3JbtEgDh+FFkRoStLf/Od6ZurPoCHaJUpp25CSJA063Mgc79bixpXCVQBk
rDTkV8GOnLFy9AzMfxsfHH4efHL87xQrxa1NCotsQnxE7U9BGQcvmZeLoCEyV0WaI8XfUuJDg/p0
EQ2vf57rF4ATgxBcNLLQ9N5OexMOyBy2sqISxBYcfTgKiIXfeN2KDmJPspYzmsnNMSk2r910P/vN
c0SGpo62t1k4zOtEkEYi/rmGkZ08Qw+nFm20pYJTUJpWCbmxAaOWL+3900kaSu8cfRgoqaw08vlE
ekOoEIXhj3qjrUi5LT8e+S1LD4wc67hk47WM2LGWTpokCDUlUQVQsneP2rsSe9PPO5citUcyssAM
jHDPhqrtVuYm+jaqg+tZlmywYBWhouYwCBwCgyQHe8XvSiSBq3cotKKP8/rK0MXK+FzmxpIgy0mf
kJJ7krW5+SJS
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
FF92Y2BScS1tYCbOJ6nl/yrS9tO5nLdkcinIUmduQUlX/rEFHoa3Ivyk0aB+kXloe21LQE4kGkQ6
Q9+cOvbtZsLXojH8eCz5LSxZZmj1OY0HgImQvBdW/AXKvPSh/8qp2AkQS6z06aDmakr4JM27sgw4
e8FcV4tuRcqkGs7bb5nTeggXj+gCM8w1pZjupaF2huj2/7utBwg2caonPL9QnFqNhJnw1y8cEijm
U2tA1t1pCHmc/cfMmTL1KVw5knK/j+GUCQdryhHqwEoaWgcU/WsJ66DlhJyiBG8LqQzPrvznCBbb
LaJ3ZRAbBz91jljSVrMpulWLCnotPmY5QRPBNQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
cqAgpvQThUsKP1YQSQ4a4I/shkrWufEhsDBDReUcDIwQgy0J3zK8Xf8BMFoFrewCsS2KNDRzQ+ER
jCDGccgdbKH/8jqChdozG61idZWa0ns7506SogoQlXjlqxzJaYEQMyNxDX7Ycmqi2PkN9cXJyFzV
5txS0QofbL3mzPtdA044rsuP1fkQj0yHft0ysK4zktjTKWnJPMDoc1p9qdrOCvbt1ZBLB18dsflT
y4tm2j7ie4QPZbNefa8AuI4j7gxnCkSCkqJB+CSn4ks4ndlDn/a3c79q59d4UozEclqodJLD4obY
Qe0wLjtJvGaBIVSj8HG9RNO8kRI3GFa3bHt0Iw==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=36576)
`pragma protect data_block
hIBljakRVoa7TrnQ7xe+CBt5tIr3koqyiE6OB8IqPuzZQ1gIn66lrZADcARxG0OLdzhb/XUNJeR0
Dh2vDmsb2cqe59Ozi7cga9PrLeyEQe+W/qJ/MuXtl7j67XtTkOJJUWL5deeXKL1VVtt4OefpB31R
BKfAqbgayqDcdhzDQgu7K85EaaQ5BJT7Rd2N7HDzrKg/heAUwsTys5FxPaHZjvNDbo+tCVpGAqLx
gjydAH+6K4tYsA69hfNjkaHwVOFUgUxpz8h/cb7TfNBWZshvzxSbftPyKXrJBafFM6GFY47OgrPy
gTyvDpmuCnFbIdqQ5nBQzXh7QO+PkoLbt+++iMN3m+T2iAMOxqWGQF7o3LqWoqb7nVOiPhvSJaca
iBwkPLpUSIB2C9uJpZzbJN9ea4oYiE+qXP3mAwCNUuCaJJt0EwGlX7acWfVwSIvu9nohGCyoMtiZ
ZXzTfJ+JaAAMUggEbVdqdZ07VycNilLUKNDodZsCZvj4n6XF3kXxY+MZgbbb57nYCTmEObik/IdO
njejVEgmx6HiTzJhYf9rpegSAXSSgCzqc6bM15Wu5fVXWOndtTEGFXFFif84xhjlWFVqeCOTMen1
8NFt0brFGbhifLO0DGgPg2LD1DdyOUzkyPUSX/wXfu4FapT1ViAMOSBxf3zADajj+Vg5vvODHaOa
jWTbFUK5n2g4m4IpcCALuEC7mwyW/Jk8QnssyAScEDDFCTP4x/dC2tBSEUV61KjFIvLOcz6n8MDn
+sVYBH0ytxYxP90h+CCcYI/2ETaveBHFEMtXyG62zEykq3LMAu1odHrMvW5rMcMSx4wW/Yb5iTv+
ydGyjCYG0Zk43ztUqmQLgiZ+sS5vddiMJC5GVim/g+t8onec9/T2IBNgzxICELqUZA7zCxdO0JfA
ZVrAmXlVSCpn2To1Fz9BCbP4/aP83kt+Y/EYm7H5BNh+apAKwG50Q5BxUaxcC1gInuZMuc92SavU
G2Gyb21ciyy6fWLdA4wmtTZC8DVNjQ9t/9hr0Wd96CUyHNrpEVrZHltjNl8623lquWhktJVkH6Wb
z+JnkpdB6TShbidr85iFMNwE4VLf+qs51jOeCUTZ2/KheFCf51GIjbnIEFIn0uy7UjABwIOr2jlx
WvyrBIYrFL/KrxiKy9Nki+HAbKbiWjxC76taGek7rURX0ROijzfiq9voHk21RR7GmWmXwn19uP94
V+Ixz5D3Rz6HtbO2Ct18C7Tm2XJLF5EZxrIALWWdww777N72cl7Rd60PKO/PRQgrc3Abzw8/HSZa
RU1YCCXBot1HvsKSrNPsZmccaTiT5EVeR+OpuJ/6Ujr5sHMxcLoskFNYhiDNHwktl8IgT4FpoUVr
zH2lcNprr5aFydWTGb1Rr2Cig/j1ivmRLmjf2ZBzXxwmGdoA1sI4mn/OAGsyaWG09dlZSr3Ur2CY
ssYJ3Z41WWiNeRtSvMdmna3gvBB0DGiZPX3E2l9jCUCN9lJxmRmMnWS95ify2gbHX1skhMLgHvaR
NOraaFIesu4uObkAgHMMk9zVToXrb/+QsccDL095RLxdhWjdNUoNFMdTVzk/vTW0Npqm/WjFBAO8
uvo6T1wcZSUvuigkhOAYppUxnYcohxS1oUGy1slYYfeLSKJnAz3Cw+hFomDGLuHmWRMSCSwM0WPd
A9Mlbsncz0LD34G6OhxK3lCiByu99DEy+3YXfcDhkQ4G2ngxrS49CC6IKNO8vgf+aWV9yfS3vjXL
UxEsQSCkkYc7JmWiW81ybCS/PUYdLxRFMP4vv2/ystXUfWdTgWSR4tFA6bpj6QXA2rYhhN51LKTm
6QLbk19C+dh87kiPFFfz3QycUA4nh7NK42AfwgK1YCCvCznLBQINFpBYVHV2wD+PS7JzyCNcAru0
GOrCWBj3PkhhKew1N4hS0dmILHyagz+dExfV5RQZeMgiZWkhj1QHmf7hRzzBTJzbek1GMtGczOTH
Gck+8l42539x5ixREiJMM1dCGXNXyeuW2aj8UVjaX10ShEWDmXI4wpDVvIsDAH+54Bv/mqEZyBA+
zozLZ8GEBkbwfzJKRO8Wt8+bFrzv324CEto6Kn4CFeXdeaANPYhkoVuzpNKxhaoBheJ3h7/izTcN
YQ0YVbLXrTNJO+owqgdhNLthVeNoyawMSO1V5gxdUv4s4yVIDXktkxODQqkeZK1wNRsQLhywtLym
jW/XsSnz2yFFK/ajFvTMUbpEWupCNi/NqXPE95qJ+vYDl7SLi3eAXO+nbAx3hUFn7oOwH9gejccp
lNUISH0NHi9d65R+LiEbVx9uFYq8BdNeK/tCQqpxFqomgbaZr2NM2HUanRdKY9EqkTiLU1c8LVOp
7EMoF4Xbbakk++AHUGkoxZz73krtrkMftT69+E51RDZ76zCKs8+mIGjkg2ofr+4FFl9alYWXEGf2
J0ZFOAFyaU2uFFrsZWMJbVaQGLbF96vu3P/lQ5Aar1/ZzrWNBb+L4tszt5L6f8Q2YqquXmHMxFp0
m+h8fZ8qVN6FRnnk4b+0/JT5ZOlaqKtYVoET2fiWKC8PVd1dTCtral6LSB/WidW5Y1q7cs5WQ3xO
yqjFKt4nlHuexNLMxsmGW/r2ul06fv2iFz+QbGeX0s0Y2aAnSGj7H2pv8nIVAHAoi1dCmjs5GFaf
pqVFzK/sgHr1tTYkl41PhZ83wp1op99vogSRr1cJ9xbDsmpB9fo017XytbweqTBbPcNoPPmSJ9Ou
pKAO1um3Yu0TSOY3+FjJuJaVnkFy5uJSfdLIE4C+WPccfeal5DbA3/zf773I4PswP+hIdDsMHLc6
nfkw5VaAeTUImm5WDfPtqlSVUj75UG0kg13XDZpEK9NC0o1uTI0FX2KaMPS7909xwad0vlxqKTg4
BQBfsJI0ZLwkUAuYF2t6fvOs+Em9jQm4YOfiqT3/2FyHyUEKhMkQ9zyAPRvTs50u1dHbq+73oY9A
Tm3r08w+Wx0AqYt8iJ7bcRBBYFYjkd7GU6UzZFIfyTtNPWrICer85eFlbR37kmBJMyyVlGGVIOjw
O4w4XjMQK/H8QXSBpE5SsM7XtkFX66F2Dr6xbreiAbUaYMGG+fmPDKCe1+qEPwb4PV5IyefU9Y3s
Oz7sX2Zh5qILVnivslBg0gcTjwNQbvvApJIisNL0BgIxEwGFcFv6PNMN5YOatiFP8kSnpShkIsW5
YeHmzFE5XdGf9r1wxbI5VtBvmR3WAYfwQK0qkNKR8PqjKyQnVmAn6VRKyxMaPWD4YLEssFdu9SVc
1ztMeYAA+CgHQ6vhGOQYjofS/H5JO/Cdrv8xZMUV2WMYSrUCIH+XsyBXThNeqx9dHCh0oh7jKjby
/5h7eL8vfyaeDUbqgJO3+JXEhmPsV6I1OawikH92P+L7pgXB2s81ndcGM87EVUzXn8Xu8friLrbr
qeFdq8RZboflLq2cscOxLcyIc3foLawGi67vKuD4pxsr5NGJ8QqUD8NpjJNXUWB2wsOsruiNyVSl
n+mJ/NCiwsIKBp7jwO6tdYxsgR9O2RM7FoexWK9ndZiYVyjucbinSFa3NZQTV2cW3pQySUvvOzpS
H/G5SQP8efa7UGQIkedFImTpoTU0l987/9KJqJZj/NiNhrgAtA/CaA/poXjx8kgbmqyuc03xSC0p
LJmkzthgSfaeltiDlQmxPahZUCEgd6YEWi5my2HZHnGD36wogRKzw9uaP+s6qXD1tGQXMYF0QDSE
/xS7xZw4PPy/zHcp30TDXqChzp6ewO4nsNi4WBnWm/PFSqsianqUek/KRDOy9lo5eRobSLabptRs
+/c3cunmfMtrr81tnTVXXgt5fZnkDTkgXA+/XtEVJvKDWB0LOkICAs8hqKe4DRdNP74Lxww3HRqb
dSCyMYnDzCdgxJIjg95EwMcFAvYz186JtmqniFFGM3L2Kg4/tw0UqhPm0Sf9kz/mdi4NoPzU84Uy
jsS+aNuvzW9ot/4OtKsgXay1J3ltM+OaWhRSIc9hXwarsziSwKA0qiZz54xFcSqY/CCtP7FnN5uY
oS+PXpzTU4nPCgR3BX5Pdh4IZdvnTmd6HXA+4MUA8ILjiMieTDPfJJMSfMFBCFHeMjnBT9VK2vF8
9huvp9HzJ66S4XSLiSzmbEpRcOnmQ2ecekxp2zlvQ+4K0nuwf/3f0WzN0LQGNnA4JEEy3nioOhlp
aNW8zq6q2IDRZ5CEQjSkMyfVZJyN1+UoNhWRLOxoshlDEdBxykK9v/fg/tGHcv2VpsTszqVWTxsM
Gd382vfGExYOCHEn64pazLKAfqzeE7TwTKmJMt2GNw8QD/HVpm499ydoWtVJeTo+I2i7CdDqpVQH
9CiDA/nfs+wwQd8CtkoA5YzuFpwN4uGPvR6vgtKu0L16FpBeiBXzKmg/Pf+Swpr+6i+F1I9wicFm
2L+NH59yTNKWzNxBV6IVOoI1B0Z9Lifc3HoMFqDsyyfDJlsivJ2HLgWjXYm+pcJcixIEgkV0deUd
aeyePcvyd2A4krBcz3JB0N6ytj47VQZtqwXVGwZ3aXTpPkpCSo4aS+w6BXCFQdgA8eO93v3Oqcft
LOKuuKex1PHmzSX2p6kHsSLJH9vR/C9UUtUrwdR6gYnh6L7OGmXZe9aPw2fr5oLyPHIEbUVKebEn
ol6msXfNcZW3xv2rZn0U9U/4GS11QZGy0eV3eWwwkigROv6mVlWqKnbV96AmNIUBdtFBZ9HwExCc
hGRz3krjx8k0+W3xH0cOgvxidfJ7UPyKp5eaWwzDdkcQcYqnfjEdQei7aHPp6z/RtbOxX91WTQdn
WlXdbuPCu0sJ+hmz9qzWK52BQVavM69YNAIvnmA6YYZNQYj3vcViqkpGpFUSupmrFDBiqaqazO/b
tk9PNg7gzf/I2n/7yuMWNFJL4o/SQ3zeF9xroiXU1oTye9L5ZAKRH+hfQRpiEwjTtUodMcpT0wDT
GO9HYnN0bQ9KPim6gXUdXH6/4FFZO4sac4mxY8Y8h35N9pwIOwUlQw/xpI3CCg1IEmwEcbULyQ8+
s0v83MbuEpIX4nxMP7lhQ/TfxvZijLw64CLaCzKDsMHYZvPzxUwd54fK5zCVxlc11RIyzT5Z4rlR
KDWShVmfS1CcE4Q11RME8UBfFI19WHcxXfuQVIFIVMV7Z64uLLnUX0wM0xEQtA0tnjruXsMXRTMW
nlrLWLvLys8oASaQTtS4XERDr3P1aTsFW7O/9orrDOoqSSCYF3+o7vCP3A1drYWKTzhEvJ7zJt+M
hECKO/qGJ2buhiZdoKFfzqzHSJBHg6Wz1KJPjqVprJRQ0afolSawyeRdSmpXHqXesX/iX1MFDb1k
t3ISDxSJpYnnJBhpzZAwMMNXHkVusDaKPCtsCbQicyUVNs/SCJRBSR/0sIjdTKygqLO+sKlLyoSR
tGn9/bd5TTL+MthwPD1Ft0flnJZF2cL5l8bgzXmAoTPr/d1jeyrGKGIin6zsciAgJfBn7t+uOo51
aLZohUYNRqA8qUbBC8wCz0MxBeD56gWtXRKbMnJ40yvWwtYxx6HxefYfBTALUm65TzAjWcfq6uRQ
rZ3n8VQskEpZq0oR4YXobcgUHEv2q4lgL9BRgvQ0w9hv7sy3DGOwRL8jDoiC32XjLM+/tyE0KLBS
UAaJt18rD3ftpf/3TO49+3yaW7oBohwV33IipHj+vaQVJq6M8Q3fG+fQm8Ff/wnQKM+YVC9JoN7R
xcWCdY0V1tQ8F1pmr4+AN7qxbH8wW9YG7x4p+pDjwo/FHI+tfM9AfX4/bpqGm3jaaHc31eAAfuvr
C+7kcHycxUR7aBD5tdsfiy36FE9HasO/Xo9q3i3JnGdfMnHKzg98h/FDumwHaAjuK78amdmWiab3
v5Ku6Trp2pB3xe67Jxv/P64pD13akg92m/wlaLmnKyT5kVID3rf9c0QXbPMgaxC3BTzvpMdds7kF
8okuk81J04WElpHaOs9FwcxpT4aO65vwEmIh+gO56FToCoQXzcbipwRP+pLjSD2ge2ghV7nA9dze
PI4j5e0iN0DUncPL0DY4C7hA5/ZJFZ14eF+Xeyxqvn//KYaxhXVrtifL3hxmazdkhRoxKsNF1S4C
pKMaYA+fdbh8D2QUtqy2Nbj7TyHoru/ZpOlAxavsvZGzjw5+qu2w4g1Paj2IE/UnucF95pUUzEQY
qq7AqVmLB5Hg4ksXz/0r5Z5yvnJGLSA5crdVFhiZar2NDSE8Gl7aRLet2dX8v0C8U7jsdwGho+aH
HCeDxcTLqaqmJmWN2R9dran1ghaFUVcstanPc3SliVSk2CTch98mYkS5FZGSVUMMzzf8Ka6nLx6I
yN6Z5BipsjE/0CVWMuLh31+h1cuNbV0PvIJdcY/vyXhuMS+D0LOVfH7Vc5wFQBRPG5dC5y+9SvbD
KUb9medCs3WKz3Ncul7gx9aoh+NZCYN/ljA+36s8kATDN8UeBpeMMEXOjVGBo+W392842ygqVPfc
cFOAujP1CDB+ElhS7euOidEKPtgfuBXTbdHws2ENa6ZmBWg+1uTsvxVyhzAJeabWYYQPQkvIfATl
4D0Z/M7gg5dldA9YM0bgh0KN87Wj/D47yDfMzY3GaQFHKwGc96yJEq4qCeygaazHyoCavu9a14cC
m8egZBUdWbbfDBvEXGaZXnaY1hrL8i8kS4P/VDojkPiwSlDs4k4v8NxWThLIL1PGB6HDiTngfKDk
4FZex5iKI7XSU4LSaFtf+jYikqmIcY50JsUUMG18Cank6sGwLe7qX8KH+tNpMlIj8iWHqQ69nbXg
t5CeeLFouS05YH975TruGiyBvgGmG5BvYnBWx2W2SJyfDnFioqm3bLtxMLHkqCngX0pMqkWpV0aS
Nu1Ou+nmKf5BJ6xh8Hjfnet5dWNBVlPCBq8ALokop9Lf7/nI3buw97TYIBYi3kWqn383HeCWcvtO
WhNcqbCnanil2zq6N3NSuAqftiSElQLfqjRaKfL7bsmOGJ2gofs7P5T9/CM+7IAv3ihUrrN9IjBp
YG9JcASt6lezOLmJQz+Jl7VWuRp6jyfp6VyUz75WzQix48xOAvDsY0vYzg91kcYV4rdtIynsBZ8f
S3qYbuw64DKt6q4zG2EbqKQkWgTpv3iTG2O/Rpf6eD4G/hVasReCI/lxCedJR6/j3FbChUiU+e7Z
+T+pOwi+LFKvk/MoXhmQdDCc9lUxHnieOETgepEHRWj9BMKK+sS8IyxRnQdMhKG6TSYYvuo2cV4i
zYtjn4Yy/1CFzijg9GvRBvmrp2EaeyPDvYWzcZ49Dbo5bylF6qkpHBm9CE8Xx447eOH7IHM6/OUN
1cO7L1tecCCx7nNKO9o9he1071Zd3Poa1alJr3bkkROS1G1XjlFixiDfLXyOd5FK2LIL3J5juXsa
F7JUnSxVrCD0TFkpnoCXFS5EPPc7TqQZ8ecR+lbKJb9hG8wrM4WqTxbkz/l5Ub0yQHfCEhDD9+VR
dgToQ2dKV62lsoa3z1+myG+XoRAAYzSDR7a5QpplvFzC3772EVs3PvJrEHqEq4fJujBAy8RCnZHZ
qNpo4AL2vn7gdOWet9UXrZR3d7X6HiyXItwqd+IJkdNybi9BbhRzz9FcXCVK73KKcWFvAKL6clYy
VHn0jNRJxVCtDvzjfsyVLJT7wLVjTACKeowvspf9v9oXG65r1Opc2dZBA67u45F32RIxwsCk59Lm
puVtY+Fk+fxowp8nPOR+U5FcFAx/rYRX9MBEdgu82wkr6nUy2ApRqGFQSEtRumblQlVynUVEKnZf
acS3Nn5P18jTtgYrCCJmoaxC7JqF4Ew+wKPenq8HJ/OFV/hLOzWjzFKzURWGfeHedHSKTe0RRqs0
KeroE6HKl/WjAQajqOZeozetRUBxUEN01lYwbnaQtBS6WzRuCC8coUZ9r3TiwH2hB1Ymn0EGjlbf
1RsNLrjcMYGi0lzRBc7XaXg5+6XfZui4JEOCaP3sMzI0SgBoGdOsmpZpaFQza+gk/fxbt4KZM3zb
puQJl9e6lioBMGUT1FX4VC2pRLVbUsgbGdufCUXcScQLcSHjh8OaoR3qCkVvTS+ov/O5Urf/F9uG
cwY6Z2lv1BRXb5Vhgbq7KKyEgyqYu4yTBiC9NmL3+lV+BaYwO0DReiG1YXvXdybRbGtJ2o2wJtLR
eT/mkruXfRZQYsyXAjNkB9/mjA1uKCUaU2f4qOTTbA+jgiuhc8L8mdqWXoDLjAFkpD3H/UoumAnR
eaWQMMt32fXfR/kxtMV7zZXVUgroSODMXrT/HWO/XNuYqu0Qde2UXnYYfp6v9jOq0yfY93sNzQIW
bAWQPq/ekB8ES5cl5GAkeX5zc31n8rzJYR1FA5uByaKTKFo0soM1MWNIAP9fP8oawx+Wh/2NOs/R
MB+OGccdLM/mmv29pqZhFSG4o4LpVLZuEc0/EaZeMq/qjpnm8Z4waOp5R18vI73gDt2/ZABdSQaY
zqZCHX7reDDX5VLiNnvbwcFCBT/9HQzvd/MFrw0muvx5C9Ggo/LuKOqkqp0jNeOKJH7h9Yr1DD51
SOPI1vQDtRLjdam1/M1fJ9aTePn3Tk0qbub6Tc3L1hfAjX2mJi6sJ/8Qv/xEaOET/SIfDFwHnyYx
cq4QmU1Wb2FFWgATZIQxQhUqAqv47mv691DfWegVaQjGlRIrZPZKd57gA84o6WYzD36BLmJTGa7/
FFYFppoSJEitAtxTwswwCbiCya9yPyp2utEOc7G8Nu7rR5u96Qap4v1btg1obRo+vRW4raH0lqzg
gvntJWlIZCi2DALh7jzJMyUHWT/pbp4yG2eRWXPDAcKkE41e3hSE0TKFbHPGKo+EKpaUvjNsvcpt
E/wTrw20grI6Uhwc7NBXtdm9iXJ3Z7joloXMi9MQFmOvokHrVibUmQu6hMOUK4zGL0sexwNczSwH
X3UqsimRitAVlOy9EiaEH5f4QVSjz2psT/NuYeF1R2uK+X2mn89h1rZZKi1NlKsqPv7xhdZMCuKF
vY2yuE5CEhsIde6w6wSZz/GqVT1pT5YMepwCG2929GLoubwm2F9fUUFDEBM3ZLWEgl8xzamuKDN8
N1tSiURryuiuCnoxQljnTNyhW+eeZycWUcN3y4qIDENMLe8ULkVMN6R10LzCGJpXNaHUK1kjfAi+
bUGeaRfizmeejvu2KUh1JInSV4yH9LZQy3J5C1FdDeweOaaZDsjTB+otj3Ii2v8Wp+oozSVf51Ev
ZwVGxJDOwsjpWv4+A8eKjAMSuXxMLrKXpZ95E8zkg2Esrhd0hT+d9YTVeq+AsP5vZmKc9gGDyebt
N1UUtgZM768TQ3Cu83aRaZ2eox+OfEoGU6e0jQ+sGvHUmOpyKrAJW4kt8MYRR2y4gGzw7rF0x5yH
8mn3lbVL9NApmhxdYGrKiUwDja5sFPy9HTwbUrvcxBvWjulZjv2YMwVEMFtPmMF8hF5eYBKM8lD9
pUPE3ULagP6THa+bxELqmCvDpEolSwPLzgVqyNuuZGYcxorKnAYbcZirWlnXXcbYJEd+unLEIuT/
X4XxI0EJ0EGxqH1HYAdZ+Z60rrkQt4vmRyQIJPjL4eT871aXLqiGFDF14mbO1pFy5DWDv0fDl+pa
YUI7Lx8THBy1nLYj/1rbAVz2fdjnxEhICwTviYQ2GgeI7K9d8zn0L25JxpT2jvKQ3Y0kEmtbEzs0
5ho/zy/joTfrE/5B4Nr0jLYkNHl0WX8i+9kDQ6PHov7JkM5PKiVdQtRrM3cN2Td5sfaPn5dsbuW3
FlKMbrxUsZjxxgg1ZzNn6sH1flKuq8Ngkn+Zkd0CAoUQqKfr39pco5VS7XiGgknsTSiykO4JIAeN
WEEJ0bJDBXgwYUmzZo1hoWxH0gyp5KPzuOEXVnb1kKOvbESRuKG/+GZT/Asf2tqV0Til/OoRf5iv
lmG7ezuNEKN2svZfRPFYqSiN1rTYb58hUPd3+Vm3TLbnR+VtAWuPGB5XyNzvOSIF2VV+AchREX69
l1NNBZaiAN38QrE4/sRs4QOjH/PXKuA1tV2sqTp9UZG7g4zAKuaQtbkecMg5HTqYqZ32OvEiZxrq
fu0oSymY6AydmmrmDhMGJtjGz6AjX0rK/2MvwMZnl6BLtoK/DafJaSX/Yx1F1LIWHCdp6Mg5FusI
tvf4RcLYOr3+OA9VwAE+5FZjoOvMvmD1qK8IjH78iFKfBL5MZPoxZAH3wmbSevwBBEF3o6ktBqI+
CGpccgBE9KEEIgdi70rHdEQR8igWQZieq0b2IOgOzmNrkKx/sL529NC5geJXV7jddbWX6r6YMyxt
kSqVKngiPfOp2dRpI5CR2kuVvVjGEZGRuCj1fypeCEAnqKFN7JZQmcZ2jut58s3oMH/3WpvNIAV1
ezBVc9/2QiahIz2Khfqe1Z9i2WMSK2DroJz2a/Z6uC5yZrCyMGBnBS2NI8FcHRkM4njG33wmwOL7
x9rJKkpNOIGYvdIhFRb3aI7XeUsCzaJs4gNRBaYxfVZUJTCtaIFFWvTdDq+BLJOzMakRsQA616F1
/yODCm2PK9bTcPy1uFKokcw8X4xgghPi7Myb2ahIzh4JmUDgmrq6Bkv28cbyklQe/mCYQhKs1eQi
EXUzsnGvBPFWybWLXXfo2iPvj7QYZbph71GdhPAWLp+Mw5jMe9EULEZf6tK5eexqb+hIFTwlJCZ4
iGTb+1AyNWy446OwA+iI5jV2tbNq7O7TEYAG0JsOtCL6myFwQkd6LABqY7o2mvkFLRuTnPUwBUxj
LVRIrunFxXBFtedHSxeEQBuI/sY3v7Igq16i0VKsN60iWYwsa/7WGi6Ej7Q92SYus3HqGIc0h9IP
KBXKPyYGOox4970WsXxK2NPY54YKUNyUfetCAWgxCjkVKFPmi9r7ADwuAIuqn/E8sIRK5kT6YmPH
Xz6qJ6ZhOkuKT/SK6i86V5GT3VeOPZtoJOzcdaaTI4kX+wjjSOk4zGHU5QUsEth18iLfl1a6dnv7
nM2GqRnVAWR42KZE/W7RYDDUgAxyrPehpc3krsgnUhZJD5Wj9ZRLU/F5Vo+o8ndin2hTyP2tjp1g
dgWOxyMI1Syq2I0fyLsh28RdnipKxIpxgAJyTYjJMxFaWMoybqz6C1zgxw3SFoAheREhgYffKBKh
DmMwOuxaJMcVjmj5+20m/HpgYBxy5GB1ceeN5HhPrelVQTSoHaaA1+U60ELvmYAJtzESbqoUbybq
Gh5YRIaAKhpw1SWzd89tTooZnVSiANMWsups3CCEcS9OR4uztCV/dpcl/SAO5kbb/uMuiWpp5UBz
oWtnuZ1U4vPfnI51sq+QQq5TAl9JxW6R5W2gQUd5wHt0JR/bQRmmroLsoNuwuDnDCDYxeQpobQCp
z/NFyK3C/kyB69MmrKXFKuMCfGXLkxNN909dbB4zeLi7F2V4HunLCzmJEIaPsEaSP6LNKjNC+szo
OU6VMouNKYjINdg9cz041lrAnneSUwXFNNYabvaZDeTDS+DxNjg/6a+LEF+y+nom0VuGyl8kQpX+
wXT7KJt97aQxFZ8lSpBJYsUo6moX1cko20R7ou3mwwJ+HePwpxt/Kde4nDHsF1+QEYXhjT+pUfTA
hBYsevnBe5edeexOD4RLHaMsgkUccWgusZ6O47ihc9XSNivlz9WLP/ww1igXqmgk1yJQSTXFWfe1
vuZg95YmyNjr+z1l5Pid3FcxliQGKZZQDhvXS5mXV8oOj7HvGUSAPphraUQ3R2RZ4/5otYRoOMKM
rsI5FoFlN6buW1oEnZHQVhsjdAGRi8Cg8aMv1kepFm0x0cHTxiQDPRVWx0/fGZKvzrrXkZiLy3Zz
VYi5Aa57KpMn3tL8Q7EZC0gJs+/0+DDbnAk7MNWrtKMPwisb1lHo1A4GxWBo4yaxj6z7bt8i2Rr6
taUZtIkFhvxw0QdVr3IY/2CkcKc6tFVc46F7ZDRDFsnWhHvzSYVJYJI+DofyQffL9zGqfmbQ7JdV
VnnoLnML46cBrR6DDtl6HR92pEgYZuw7cge/4Ya5YRlQTii8sN2qorT1+u1S4XxwqnXEAMyQTBvw
Rm6CiNaKQghINNZRHbbfeErESEocXHeNM/zWE+dfLU2vLFnO8zGwWI/2I1RgjfqzEdx+kAQ9Lu4G
4yqPlnd6LbPOD3uti/xRtpgBalUGm35V3kb37Mvxd1dzyLSUkVuiXF4saYCYQiXvhFsGw2X1YS8d
J/xxTVlzS8JRDvE/LvRkLQCvvsehNdb+fHZh3yRf1fKluVcDGNLG11c3Y3zTmBs4w4TS4Cddx/7D
aH9iDfccmCX76i4DSJw8OraLfCzYXpuPEjKQBHx5hceTug5acUg8n4ysdiSkf6H4usGEZ1ZPleAs
Ww4Bm2IGLtKkRm0UADUsFQerslVnPKXWxzZUaZ4CiNBsBmZF/w6Zidsi3LBNASPyDzIta/1oBnP4
xALVGzqF2Tf4MLXJxXVGUspSRKkOXJev2VkLCibuVBVVD4ITsMaLipKb7IwRNQns1vdsUadb+MEf
2UOQaZj2TTBFkzmPtesXHjVaAyHYMqMOhZ3gVAW3XC7sMLEIeFbC7vzPzSddom5cLd4zyJxf1Ozr
Lk9DKjCu/QEPNi7IB+aLg0vDit0rblAwRaCvBhcoZ9MVlud6sFv0Vun9+Fs59eEENUt1zrkV8b7n
K8L7jt84Y96MUO4Fx0/9/RpKw5q2sw7ZlCJ2jBuOPYLVIHMn0Z5MW2ScJDYaGCGy4Z9UMFp+9kkl
uDLaC6TonS2rms2xlIUNwpFck/fvl6Lg75pNvFxzCgnvp3DlxI+M6cIkR8YWxWndIFGng0shiYqD
ecpbfKuzp1+twwyvHO+IU72JsKrJH1v/vfbFpq1bN3/UfxWEEpk7EihHsg0+BSpiS2uUEo5biN6O
iw3FZ9A0g5tbdmyWNqZuwNS0KJuiwgV95f1U7LLxHuFTlSrdZ2sgyKhSnnKbB+eAwnqOA8hP4ZPo
EFw7Mzt4DS8qq05tZyNjJjcrbhZEEVv1e8y23Eo/QAfEy/AdnLKjiShAAC+Kr1ED+IuGhjiRQire
v88m8DWFwVJeLYKiWJMGe2DXQVthiMYv26i7FWLrUnBn/M7CUzOUXHyDzECNA/pFb86NuGDSQucr
kymlkIDOttOuMeAiQI0rYdgrBXZ9xJ6oxjw+hvMJ+IpL2tV14T7AxvwwQdKIiSQKsLzB7lxKel5w
UVt34Vd0hW0Or2HXC+TdmtxtlyIiGqC0JNsT51nHk+ml+2ipW8rlQ/SupNaTGyPoFv6UOwAv2/6P
QjlEuUJRsua5Y8lluz/YAU/SJZjeCwkgkksL5EJZaYQbjjfdlkKGLEEcDJ6n0z7+phTVECYHeY9k
X/AVThzbFyVsBA48K0eW1FsS5S1ayzsCipw1wpyr7cNoHVqd/lOe41l4RYkigSeolCK7WXdrY+tu
nSVaBqcMz74ynV69LXXdQfQ1VvjOaJL1HVeZsSNoT0+avt2RV9deyDHqmxKlYtgTfNLe6GYqTgJU
YjRA3XynWleLRXewsG5UHAVwCcs/WTQEo4wxO2WVj1+jvJCnH1sOD9bA8RPjtLkRvTS84ZdaoNPr
d6gD8+C/UBCp6b/AARVElwKkRqU0hyL/AzYhwjq28IrQSpucqrbfzUninHmNz4AaWbFoObfOkIWp
9T/YoZwE/tPYHGifY0TSHHfyZTO28594GnF4KBwQAgeLCsQfrslp6k6xFTL3/4if6nOK04KyBuDL
kfqH1m54XGUuGCUa9uPDc2JooG6m16qrAkhWLrBW4bDwIHWxIfZQ13AhSeBk6X220Wc1YLv2oegE
AfMrSz4jQOuRSu1w5CaVKc6LlQ6cbOv/ytel6LUArYWN9GlbmXYxlFkEfUU7dXdcYBz7r24fGi7B
TSIHI883TM3VajX8EWtFlvR6Ib2hgTbKeLBQjU+bzJ4FvGOSJUwJmfeRd+Mwdz6D8II70PKEGlMY
WwUNObjPYMdlxX8r6mxno30gm2me0d0UnhE7SzHvDEpq0f2KCcCcOMLXBsd9AAHOUTdTb1dVjdiV
OHThg9qBYZUMIF/PMoY/vqvy56kZ++JHyuo6s9/ugOS740jIvh+iqkPLShDxFmgo1Jtsb8kp35dv
aIOpgZ6xV9sAYCgyLBBuDDPnK/znB5L55Td64KuwdgeJcoYj18W+lokj54J6wOq/9olBAue/FJha
Qd9WFLsD7HIMKuGPyb3uDBk7mKfxtd4shX7oxm5HfAgZCaYF7oauspNDj5jdxFsF+lP+9oy4wx8j
Q++DyH9fp3oWx7bQcrlST7ynpqnMvw4x80AiEwJZ8TFStLGb7UUY5TJb6JVQRJ1H4Yn3c3dP+Bcy
9J2YLl/0XVRyAyJpn0aupsEPhDrSn37SheEhxONsSpyo4eAdrFWRZqm9zdOiPB7Omy9rwnRbdjwa
E1fhy7CHf+5hd/VAULsyW4pfPr3hP3IEq0lau7hQH03JoBopqt0P4yG0LY5QA0Ez+2eNimDuDJp2
Ma5aUVvtzAcHJWh3xn6grwqvKpx48PU+cH0J6H8eLc5NVkYwk9T6w4qB/YfHAvP6bTzkbNIXnhTy
cpJA4YaJpDgc4sBAfjSbA1SLaS/YVRDVL5TbH9pZWXb3LYTNuuef4TcyxHUplAR+3oJxJM5vLORI
h6sEz6ERoKoHQLdLs1nqpe74kf+EbP//jSrucG7KrBtCcAvgQAO7IXH8XVMk35h31P75Pask6lFw
tqSBGvRLEZRnvhnfZI68ohqjs8Ew2JLFi+CwD36fVhlM1cnMquhjAqfA8SuvfydP43XS7gYciRxU
prw5/76/RuZQLKwxoonjYrOL+77BbskrK5RfONq52XhbMkGiF2zRv54Ni7N9DDuU95oEq5q7Yq/G
rekk5Z39qjmn8zbsdXpX+d5ZgQbQ0wemUVJtHX+ItcnhU0to4cClWFvjtDhS8UHMAy+2dCGpNubU
Qmmtev8rxE6fL4GVailftcIOZ68u4MdVvl3nCh+urFQk1hj7FBUwlvMTK44RgBAH/oQGCG7C7PoL
SldNragmS1CgUk3A/StHKGf5AGH/GwG0VEbYrzlY2wd+MKvLyjJviE5JsUAaLhfLghXvkyNorYJC
ED6yaOfPyqcMxvOvs8RHgI5jItf8SrZJplbTj5d9ljzk2+icFzwB9cxweosO7AMHI1ceZMPoC1P0
t0wRyaZs1/5PftP9vAhrcT4n0NhHKGiem068Sz4p2VDL35LB+nmfq73evRtEXD3h/bfZaZI0QbXi
KfZfSPqKzCUza7TUkqjHBWjPtZocejX9TDdrN804CvKzf49zsdh7ga5b7iGKLZU4obXoT0uqsfJn
/f8KoUYm1uE2ali9v+gzaM7XqqMsudwzZ49NkN2NA6CAj1waNaTSr3E20j9+rl6v7WfxU1AMb3yQ
4cn7zk0qXD4bARphZJFUyZ/GwiItZn+/fK5+K61VWX6cjBdqNSltOuPfw1wTodEUeMTTwWWnw4cx
xMOQSKp7h6+ilLyc/lmxAi3HNr2BpO6kt/2o4ncHTpOTe4kHRkPwSItxXUPNWrFUoQDXWyr9r9es
JeqN2OMO0k0mvpptc6dblL42tmJp3bwdHWIGWyJJOwRZA7aTgC1pDw/rxqldWYsD2Aeq/I5qr1So
MteIycZ6akQoU8IygmHcffkTfYoJf0aBgiJSatvjNy/fNZU52oHU1dnSlJU2QQJHg5a/70rhiWBs
pZx1WswuAQH8SK+hTENLLfUCLJXk3CmbWn7divLbI5o4ahlMunM7awSlupTKWfLo/k7KD4PKu/aE
9Du3qu8R7MDAaGDA1hvnrjdXMLOzvymgktfYbeBST/ZZNmsFOkOtO6QGqm5dsuqFhvNb8JfNNtbZ
vH5kO7Frl3XHfYfLP3fOl5V/AxqFrLuxYUQJ2jfGqGOZ3dil5RpGjyR/k0ldNqpy880BlHG96siI
Pqsz0JL5ZSiRs4R8dR+mtCGoBKbYr3g1YfsPzSUOfKjprgiEKZi3vMg0O/phTZdXpBzkmW+ET6mD
2GwD1cTmPtn14csXXXsQj5kXiJESnp/DM2lUlZFiGEdsYfUBtmuB3hD6bLv58StzJBYcwA0cv1Gg
/q4zU1TiJmyplqEhSghBdzVoji8vat8pxki0ie07LA3dQ0GuAYuRFfeIbiEjW6NAsR3T4838r+EY
KD8kmT7qmlXK1GJmR+EZR2319iMMG1lDIcl6ZEmmy8n3WytiwYp4qOeGu7LImzmIgtdmQ6EcRxkz
5T7Qio/s1PKf7lJL7qWUHSnmy4YnafxgudTB+02xQf6rAG40CojEsoT4fThyvumUMCzcguv70xUs
JUm3wC+3YkHvAR+gtRt3UO7jtfNQjcqmi+OydyK8piWTesDrQNKMcKLPi1JdfvhCvRM5VKt1c4Q0
whpyawJeXJVDkBMFoYmIsZ6DC0f7klv3h22BzUGnhJp9Z2sLFa+tbv0MbAoy+yYU3tQHSPpiJAxs
dXvyd2i7hqLFwi6NxSrGypodSHU5qYPkdEyoiDxWOZleJNK212m1yw7lSEFUfwKxn9mrOSvQE+g+
g0FTXrf9dPG1fR4fQI7rNaw9lcYyYNwlk8MpYGLTZXsTWOprOK/lcumWHZ9YMAMBM2WQBVUj/4Jv
5Mk9XndW/TaU2B+kFKHdSF6ZfUPhA0F9Q/Z09dGgf3PVacks2sVHQleeCNONdhYx1m3+qbXCQyw/
CkAdNt4OEAQNH5L2DyhMsmdnj4DjCKBBm9h1tCZ0IHZfuiutx+saMy+xbu+M5csM72glGNL46D/i
LDFvk0sMS4fH62e1vGEM3rM+nCr+8XrsLMRWcaMCgi3C4ON5KyJmwQ72hxCmuHgz1NvaaL4P0sfw
jDElY5f0v5EKuO0L8mVDVFmsWiYAO9Tnj7SK7s5pQXLMioF7CPyvhxeI0hGLi/orAa8fUMF5zXOW
dHpQQQqVXs5PXD+M9ZdnEY6gB6was9LFtuV4AeybQ11quxh+cHq8H0VYiT6utoYpTriqxypRbUFw
+kh4rTo+NqQhE5oEjKheD9mCJoGSGjvQ9zmM1krFX/RE/G+YhTl7UkTiABZy/6xdaPFtn8TOT64P
K9SuaihR2N5CmYMbAWGuXqwDZBeydXeOmw2lJhl0vWnybuR9bbGK13i1FPjgkeRrm2gelbx0UrmU
a2p36XtXwkcT899aoS94cQNHJpRLLUQCWzw1CrVW3YWdJPsV01EnJ0F1AG+Rakt8yo4jQwhitzkD
riaA2ulEI6m3Of1K1e40ND81KV/Rmrv4uRSJpPjoe4m9zRTslDNJYvS6N56n1CjsZ4nztWfXu1lr
GJCVKY5a6bG6rOPUorsJVbWtkCgO4SHMhR+NrLsomVwC2kyLuEqdneQoPPh7x4RA/8AVuQetDc8j
aBx7mtm0GWqF8fKz4wyk/vTtzFKot5XhMTTNYzoe8MeKa2VJet6lntR1w57l0xD6jL660f4V+TcY
XE4bkcDDR0GmHnsZO53S8wCeihLETPtFokWXzNK/09xz4fOVmT9ijt49SDwTJPfxf2CRtaV7Q/Ln
5fdGZ27TTgg7vOBT9kR9HaktesJaKW9EegwN4iaWjQ4x6dzsbMHmT+aymY7p3yjawYTUePqGmWLI
AKW58a0enLDbO4DbKxxGleNYXRH1QfKpuV3J9mGqqtIv1wpnd/UKDiXla5Daf11V+gkPk71/CYL0
2g0oFkr8YIzis6wXb6bEx+UoQm2FB/EM1V6wlx9dOZnGZHjE3iMwi6oeN/jqrqxr2slCHP8Nmzvo
aB/381IfG4vX66DnuCule+oHP5SnYCUL+KEbiM1NEfN7r6cUuu+Izh58uc0IQY/Ie+jGUjsSpyn7
ArCsgXg/Qc6pjgrHVd+ighJqO8abw94Egu9AGdv+i1TiOs60FGu925ecmO1v5a2+uK4HxSbkmCnq
6IGsNvBiZyKmbu7btz3vAs0nWpD2phxbT32i5xPfGznCEYeWe8ehee2U1EgSpJtJ/LncgaB56PVL
iDliVmWvG+2f2IBxSbUQoQA09Xu4Zy3lfQRxBXhsM4oVSULaAVeF/HRw+fxdYCTZc0I7ec6ZbftL
ml2D3vCI/PUgmY8fFaK4FrB8aOg7lhFQBj7iSSMV3ldSJFkKnbahW90YDNa9fh3/cMy1x0guLZSc
zAy0TfGkb0xu0Ij47eDrJ/fm9hB2ldzUN8zOb0bydEDt8Q2j4+koJQNsgEJ2rSZALLtLMsz9j76f
/Sf0KZzPm0sGH9fDGXuKteirgE8LyD2SXW9WIM89VuRINEddHaNJavQmef617AvIEWxNaoglVHTV
G9qUhQENXn5sOm28mWLV1CLmajzN+/k/i9HzxzJelJiudDvKalth02Dm3NWZcX1KSyB94ZqrItlg
atUgTdOBgbxI6/lbrgq0L7azX9OBgbvn7URD/eP4/lc9yHAMhM/+U4kRwTD9xWSpyglYAZjJoAiH
AMvhktA7GBrcgyoAulFiRszXJ065ORMEj3HviftO9dvleyWH03CF63Dyhjg2Zq3aC3TSjIQOsMs2
d8yW809uHlFlmT3RrePHG7/jc+z6BuYAkdJXQjugVbOhDC4mqEcKZMsDXdLzxFmF7FScvIN0kXM3
I5vwYZzHqocaI62QLWMsivGQ52h6W29ZurI1i4HDMdtOVWaR96tU2TiDv7JavFUGxtmfh8gHPm2u
/4Kw6GW0E50X9kgiJjpB+uLgzWMnnfyzR8JElWkGt2S+kr66pgEI43jyIqzalAVuRBpTUl/dwd38
BJRYuZJSXZx3Wyqt/5jCG58Gt28NSSoInCvAAZ1byAIFU6OXKMyiCOc7SxNX+/kccki+1KKJMMwg
Y9DfQpB/wglXC5ItzmykS+jRh7xsNWaVAviTwZ/BEbFJdIEKyqc0Scbct9ZepMKW5DNH0XX4Dyf/
D5tboi45bCRl+Rz0J3AuKQo6aTIjlvph2yhGO3DD58Suv0FBoiNnWbzoeRe/gLzZkRAEhaoWdLTv
m9gRz0aOMeAB1TgCyTB0a04auGM9E1rHqP358qGPdOL9BEONgAb0TlwpXpgprFTk/whVrc4fpSO7
c1Q6i7fC//SyCVbOqNtYySX118EvsRYxq5oZhF56GC40qIHyrrZeBK90arqUq1mdZIH6HF2qiNEB
CzkKAYcIXBqhwhehPwKnrYd0TBRtSUvILZgVaxDoOLbjBXA9qLCboeUjxQQtGwZhIZ5RcO8/5toi
w/O+Nm9LhW3YfkVoX2d06pHdnQ+uhxwCZXKjjTVLAc9VqJqjrkhzV6G2fpgCIcugu6C9AKK/gbM9
eC5wunOKFckb0gUTdv17QYm9xtHjPFNkanjJ6uGRPMkqg5bPlIABwKRCxZgbKZH9C0eYrFN3R2ea
2dCu9CLDAlm6kDGblnj3MCFu8/xPMVNAmEaUCv7hDVOF5BEyB1AMqWV7A6l5fAO3v2YhGYsHkr77
l2W5WePnEBjHPb7PNlp0+Vci1JL4kaL8WYOs6Hq49nBvpfUoAKLbj68vytZbCc2LwFsxDRhzEAPc
s0FmFTolNTqD8Gusl5xAUhYYJCoF+6s6BIUcMBpHiIJaCkumt0W5oR4oxgSibNomI/MWu5Z7B05D
jLNv1yA9RMAppty8O+IUqBQZH0fw46hXybgiYexgq6x+u6pvMlpXbXbVQdkA1qFymIy7e+e7Ys97
64FJgRHoiTMayDsbK51sizt14fkIXIAY4B6cdNUDckcihIhzy1q4xjQ90fS2Mirao2lOP39FYkYO
A8ycmT7UOt1fPI2e8Ky/1fIreNzAAm9ao+X6CAPyPfDcyxtCj8MFa7h4KQB9bVPSkjFNt77Fte1F
Q3o3UoPYhApEz8KnCwvpnR1/1daSqetEMRBZXrZPSY/4ntz6zXe596fEeucWy/RlkriLwP/NQyaf
O6MwaSIUoMWGm8gmtfPRpjP8+gMBFPb/PXO6NhDwO3Dj9gesxWnkmnd6/P3fl83KIA6U6jT64Vug
380F30vQefvJ9Yz5/KID/JKYpod14jQN93mtqRmer0esIyFhzlMpI5rySO+caC9GRBnhjUuJrQeY
kgLkzDn21Yi9OJkNT7WPzID2kdSYRiobLzKufGqi/EAeeaVHlu9wrX4+tiadLEGRv++MNC5VdnW9
TLkq1YdEjR4WIVoNd4I1JPd9pAIAAHcpcwWnGi9d747ntOBy7wektzpsMwqCmm+Rl7HwwYvmya/z
sqVQSkLQg24GOOzZ2l0Va6DwgLnq4zPcS5htkHipQinRdLVErM+k8TSXcIh+ycUhBcYNcrjLfWY+
GLPJJIZFYf0rzRLBohc8/TLNREVPfkUOMTAUIyFzmqXdRAlzU8e/m2CpWd4mugZvVqkF0gChzjKF
VWPQzf7YxjNv+eE8nZg0tio2ANLRNopnxhLVmB1dBdoc5UqzqrG+OWDB6C9Dgd4MGXxoslesTDBa
XaMaWmvFSC/uhzbXCtWYjBEqtPSnoBGGTRt2NQAVwWu73k068QTnTe5moE+OV6YVRQk1DsyCt/aO
r++ImH2tFLz2RxeqkrQFPWD+F90DF3DnFRRWLoIsDJz75/HfohkvxIge11ph1uWczMSpCCU14Cbn
iV/wW7Pa9IngLo5GZ66tob+xiN84Xrn3Jsk+bffj0jBvmkKCpEUz5jiuX0bNb6dwzHKtsTb4nZ1r
Fv4gGvgp+UVM2yrI/Qw026LnGLaY1G3IO1YyZ5G65eLJ5rXxjrFncwEl6yxxAinrG+O6scOT4P13
3AisVbu7zlSBSmXdMYYHutE8dphYzlGcjt4pOWBL8O/BK7D9CMhFAoKuX0zSDvESe01e0zGiuGSX
xrZJgMeuLKbFb7gNLTr4vhlTCRM4A2wFqxw2EW6kO3n+84ZE+gJfmD19XKj1mZJpbPxmZi2UqN/E
E507iQ7x5HYIgqBEQtKPwTNq6gUVd3P//LJrnRIrb4NuLQEe2lIM7at4x9yhcHKZvOSZdaYq2uZh
fZb2SmpAlrj35VOMtsF90UmDcd/gUUoAPpCyvhNH8Ec6ByXsySngekc4Jh09Vk6oz+SNUR6dyBT/
VJEz3/zipKLDOkJPu417RROYOnVDB0tnvx+Q7TlJuyv71qc3Fv155KSgAbmmnsb6s6GhBpOHNTbj
CNqNVCfFcQ8dnTVM5BVBirNQf7RDIaZt1U9dgfj+sv1qHWUawbShGYcDAi4EoprrTZTaJ+cshC/B
r9Cz4Y/VBMv09+FEhK0EC3B6SclpDNECm26yTekVotrL/e9rgYhF+l8tAzNQ9Ce5tP7xsbAjPJyc
VlhnvFdSVBlII8FwLqAICXDWMIaDj2pKA2Y2+oYQXfIPcfuyyYogxrU+S1clilEK/jXnGhezttzP
B/4/MgRPVwzcv0wryiPXBU6upIiOeAlvIpNVUtUKNjkY9IvsAtvfi/ZjHL5XC/NSfY5NWQL9KY2u
vHvvZNUD/1t/8hUuO9g7pN2nHSO5U7n/pFu3QzsLWsFWgIrq4O/sdV2n5haQV493ncHFCkh1QW0K
VwhI66+CkLPjpKE6C3Bmf44D6KRcC6/c/OP6zNRWQ9Cy9ljZmboNQFQdtZvDpk0X083BMRIDq2+h
6qY1MUw3stRnFVtb2LhcKhNlRLUi6twkxoXejaA23IT6o2hoCKNxXiR7zeI7u/QKpgQ+piVv7Pdj
DF+D9CgKQDzisi3dz9xNAxN0x7D0MQxIWviwf02ojZTxyt4AuWHyBZgACemH+eXVxIkxcD8Uq9M/
IClNc3b4fXvpsV/0iKvsVFQ6XtKdtZY3oUFvf9go4ic+EOwgLgZhyOYW+PAH80P9QbarYVBYXpO4
2CcHEXM2isM7s4IlIM/r6D05A3G6iEFDr9O5huScaEaYGwCj2kgSJk2fdpo2DArqrVjxkTg7+jHh
sHLsJBNWAP0XdHnbc20mMm05Zx76MR5jB1PQYhgSjEmisA8h4UhdVke/uNVh7cBza0C5yy1Yv/k5
FEfYU+NiarMFNriSz3t/disCsBr8aHXemCLRBh6qDcbHvfPQz7OwzhTcuQvM0HSL96tXWjkg3faF
YPVVte0I1uyBcCiOHYA2wk/RYH0cADyaPtr4yRIcUxmlEIjGWHesZYuinyNGYBIMNBRlgXFcCyRF
KowsbgkKNXAVg/mU3i0RXEpi8E/b7sxkLiakk3KuwUdpsQcqEuqoIxGsNvImKUUsq1A/BlfdoICW
Pjic8YJ0SZRlsvH4557aIAK89rSzhsIJLjmex7YpxeymfwAa+DhUza0m0nqQzCxIKTYylJ0VWh+H
Qkvl7eu4+auTy2xFT4mTLXO0M7gRPFNyh8kWbR0umGV8vSCJnNKgxQ+qdQvj02IdlvWCKcsCtJZd
Hwji+j613jD7umgYOhxcdshH+IaeBMKOXK8Ek0z1IV66HOj7k0r9K/b/Ze9X4S4beb6mVpoOHczm
G54hMpr10SbfqgbOBceBQhZpbNi0eU9/ky6OAoE9F1dZ1wV1cUv/XfGAJnbuMR3bpZWDqcYo6nWg
rG4r7YAs6quobom0Xv63tSIGmSp6X4mqxLQxwXCCaP/+Qo2ffGR0g4F1Nq3XVlQAbtDPKisue0Z8
ib6hLLl53Ruzu4lsHOcnUT0y+7J7N0taL256pUsTaSZO7tPkE/k50vU5hNMPeg3e/fZrBKhuTpmx
71PUgSwtwt5rfE1+W5uWu8W+BQLO+7uQHbcrR5ME6waNL4GdATHouQjKe0xqUhy8v6iBoHbLrTJg
w3nknAQeeocLU2cafLe2B5kZ1l/uIiSnYZjf/qgUHHDG93Kfb+jtOnu48zquUylE2uycTAXUAgZB
edZRIc78XGisvZJ/8uLk6WVP9s4Z83N6i6aBvPVCgSO71FxM5grfmWU+GfRWDAnZuU+c3Ek+BCD9
CCaVB7HXqA81Ez6wAlW7IU9xqKeY2BWStbL/Zd+ELobN1o3s4GFzLvM9e3lK8MGfXls2O+C2af6M
5fNUzhFjnk32VIBzZWMM9oij5cvcUgLKaAgtAX4KNxnk0IspGL9lIYQF5yMIj9abE5c8hbRyryIR
xUYLzwFeWzhOmUX5PZQTZ238Shn2AO51Eix4owGmo/G0z6MhpFJLkE4Iv4IOeuAGGbaKa8ryokbX
U9VaPczc2qVFPb/LqLHe2vF+rULC8fF0EK+3t26sdHEc0JQqCC6o/3VNl/zBjv3nOKJGEktOKOJI
rqU32tQFbx62Uv2HshPUfRCUo47baWGcPNOfhOm21nAxRF3eUBuO450dbq+JkzWuOdEye01AeRG0
gpZ4iwFlQLdvGY27p1BH//KujXn+PQU6ll4ElYaE9rg0fFYx1kFDexuInt5XLwODClNXX8lTi5Ph
0TLFRTfva/3ZfEy0NOP5AjDKPxM47GVCCH7Pxw8jh8cnShuUOMcWeyCY4NQd/uTmDfarY/hnUjFF
x/CNqy+45BLrmQ4iyWZTFx2f8Mp5ktG0oH7NRsy4JSEb2CYXczzrt6TdHgZ9E+YFojsNTIa9rrr3
kiTyjYJW2DwJC/rLU7qV6JnVcVKKWkKQT5dTZCRmXod2jrtef2xpKjwuZwRXx3yYAz8qtTUsBxnZ
ZGlIgAqog7OSjd6j6i90hf4EKsIf2ZvxtSD5WIygpuE0RG26vp6f6gtvIre8gRVugz7QU95P9ZhG
zJBVhcaHvaymTOBq6573Z59zeIg0XefeLUCIItcVKSioWl/vHUDTGQZzDlEJ1MD30axciIA15MCn
/krQq7LhkJhv7sNuobjYEEXTe1bOyopa4D0ghOoCsNn8nP8jyttiMTVP+rvpqBxCeqKjV06OnBZB
BjDUnHmu11FmpS+6cv32evOvNEuvMgj/oT8aDex+F0RpkNuU+OrBbwYyMS18wfwAcpDs1AFVAqis
cznXJh2o6OoTMKnEeIex7Tm26AJ2PW2ZXysnJxkw/blW99/xygWwW2OfJaKEj8yqIo966ELWu22j
gyJT1Tj3C+YPMd8UX0qSH6PzOz1k+WAZtEq0pBZsrRljAwMdvWf/Rs8TjTaipi4ZIJGHNDqSa24A
Nd8pSFxnlbEnbUfcwv5Jd43zdfCSmb4W/EW7l6EHttln+gfZWrl21aW5o9YiXVKJaVTeK0Xd9a30
PZXiyGwVblbaiSLC3fzdBBXjf8FNynfAHtqwdGH9vQYyLyH459R1C9R4vy/XLhdUJJpzeLpwfBSt
BygXUv2eQUr9+B0peXrPeYBtFqIJj+JLgKlfCy9s1RRCtWYgHpyFHGUefqO54qdYMg5dzwbHW3u4
XTJLuZIdOzSZaM4236N69xhKGfO0q2W3rRz9XlKKjfNDmbVoNw7raY1nsXf9A7hfCQS4NYVf3bDz
Qh/wCmnI6fwMD5YsfO3zLOA7rMtfVg1HpScb/9jwFyErBlyLIo71y66AroNNFaaQmSh1aZtij0X7
fQFuhU1f794Q2DgyvBMEpb85g0zQXe4ffwgTeNHbjXTEnak3RR+GGzIOUVGZa5qxNfrT4kUy9dHx
J+e86Y30d5c2K8/RVAWxGTcEWr22M4Nahwd1favT0OtoijohefGvYy7noWrDd1Y9fLp1MO0/LWxN
RgcHZ4nDIDFUp/pLh03dvZjJXTSfrrceUsyi8qhH5IGk3WsvcCUarE31fP87WrhnW00UlWknt/C3
ayTC4Bd97sx1uukTt89j2sTsWElV2/sy3n5InjrO0di9Yoif4++palSA3Qe1gZBY8nvDiYr6wZnu
56rByhZU6DUp7qa/4tlpn0F3l9pAoJhYkm3b9UXoO74MMuUpL8OW2vj6R4wNv2W3lkPXaF+fKUJr
339UsF433Tb3+pOrUvxtsDyJaDZA2+USlQb0M5y0IOnHY5wcspS9rAsRPKCwYo6ixhj/aoM1aTnt
a5L5mYxZn1O2/Qjd5V5Fqd9KuBO7KhEMPbvQ99pZQGX6wK2Q1NNMudRyeMDWbjgRe7LLPR5GCSxV
XZMIAjUZxD7vIkDcJ5yOolyqUVwFpDI5L/OWq2NsrY/Mh0Q88e2Uty0Y+9ny76iDBxTLmd9lt6n3
VhL1c1eEnQtZCddSewamzc/aQSJfEgkUXL3LOQDqpHugYcPea4I4gHQ8gnCBJ0Zgq6lwy3uroCiu
O3vfBhh4E62QMS1pWUI4Ymth0tNn3DhYwYvxXoLTQAQbRDMeO7BAu/cJ2PYHC967uzNcOs2QkYAK
m5joazmB7gmoZgc6R8Zc/3Jl4l2CBchP+2FlAMB1oP9vWSk2H+QDrFVTeVcQ/3bnJxB7SVmCgJeL
MoS0u9ROQuBEULnbJZ0qXGcqvoaSppKU0GjNPpDzBPXKpQdg831iGxf99objimqAEo1eS5uviP8U
sIBVMb3ceotXBuXNMoBNkOeLElIvEQRfzP8RfarcKd0AnpLxwupt+IKyVEDTuhA2LsFSWtWL8t08
agKZ8TOgYLmYWXOeq5M2kSgyuOm/Jebkp+hzSHcHHfNDpO+8LD9feq1Qw4WxJosdBSdkTBwXKBke
1GRcs8sBTe4uHa7+ORhLd5aXMz9UhA2A50Zwo4cIQWyj6UbAgaWOWQEymQn6jUBdkcBjR4AmN1Yc
64t07ASoF7fst6A9h2J25p0CiFo8n4PmZAH/ITv8z9WuB0wUVtwY3mSHtswsGsB19I2YQXRw587v
3N7L2J9+xUqDUQ6/fBggC4+BiMp9j2dfjC05/ntIuGgVPqhqQVmIGejp5aZ/a27vfhRoFIGMRFrw
WAAS8dgVQVqZCMuqqQZpN3rn0wbBOeN1eAVeLCawKcJfS6MvcaKKIUb8S+xjVuKFd34nYGD6564y
kOg4GypMOdNj2u7YIYu8Abz3PqPPnGLOm4suq9VvJD4sYfacrbPwVyD9bytRk8hSs/2FFla+xnDA
yOTHTMWU8dptWRqWAMlZk/SJmTZfPSUW0u7NaVGFs6wEIWhMsC4sSnAD5/uANtUHrslAb16TJ5ag
nZl37iWBx1i/LGBz62iKd/65g6Xhgc9hwFu6KW88kptgWG623568ZurNuVHx54phrgcFYykqbZaF
5pY2PA8ac5b7vCxCMgZo5zpy4N/xyVmRU1qwsqFTMGT8F5E3FESgOYbXoEcs07Y30IXX07a1V4/p
+B8OwFFOIQrFvGd1KPfoZ9biVHozYp1gF8X8trzsBrJZTF9aV6ONHpsb0L7ZZ+qMOB3J3T9Vh2LA
fjgOd0DMvRGQgYMA9Cg9OhkfJH8oqCNzHZnBvHwSj/pPirSEutge4id2ksBTJN249UGzWQD6W6O4
VwFmKiAkqjSutu/+Qas3N5R9+21F3ZRuEAtwmBGE5DYZyt08Ctgk0rJmU21OU+9O/8f+oPBd/i/J
J72JmhZOQa7SWvJDlXL8qIg1NaVcGDJM/NNJEHckTjUlKniWgUewV4mDUNB/Lr3a4itYtIkVanKJ
vGaoFw36nNotI8zqWrV/cb8TpHNxvP3I6+lcrOmcgXE2kbEzKcqDZI0Uzm0OcMeBSnCNnvA6GWsb
PgqZIuQU35pwAcQzaWjxqO+oPvWDXF/l5oK5UEIgNW/GAoaOugdXgxHy0JGDYZ3eTks3fopiaOfq
Kdbfto6J2m8W6Vu7ULsbjAmzAj0+EwCprcI8IH16WBSlQ8Wbh2nY9LZevyI7CpD9UPwOvuGZejJw
g7PbHun9EXxPaoAzZICOJheDqD+kSQTcF+cln5qDf+JEaglHBK57pGb8FoJUObv46ntumlFz75DF
FF/KYm2Rci1JZQeKDGwU/VDK0ZlchPa/yfocez8xZJNur5ioyJtfdWeNRtqemk+/eldI7pkqjvKt
ZW2IO8DoqwsaEU63FRGUByP9JvI5cIyGQUd3X77bZPepsLIv+Y4gWdyu3NW7ERhD8V1sL52593Gy
d+3W3vjCCqddA1K/1tmh5HmjLRRr8xoaDGwVJYfX0QShzab8XX5W3kKVzLr1o6sEw7Ucb2xn1K0k
OEamlditQZ01tkocvronDOIhtbwFmQn9lLza2dCQD/V21wBLCzce/pTVBlyGdnMLeenxM7svbLsi
E5TxJ9oWD5TaysrSxej9qmfLTwuOJIcM4ty949YmcgeUAt8qYdoX4BV2x+Fx+S78rbYZRSu0Lxe7
ghgTV55rXNUosdKjhr7vYE3OrPIG0XskkcP5QM3xwN9iczKgHe5r/EqPmD+Ik+lhed9IK2Tp092I
3P/JU+B6Iw02qL2fUXfgNjboY3t+z5Q9IjBki8FL+tK/oCe9FWwqfN4624TiEc/i3/htFyNoYyTm
PoCGWZKIDZa9UHBDu6UBJV4web+c4oJoTSwjbyDISh/CwuU9OS/bA6hbsMGNx7xhBsR4lRmV6UlJ
SLMlc/CCLaRSDVeEoeQOBQri4sKWg90p2hFt5u73p7VhY71D/J77obyZFfJF7eLVhlXOdKSnVcdJ
XNREaOoMEh+ZWNHTVv/EEo7v5koNCTQmGSHl1glOxG/JyPIlw9Ufhcv3cYFUUBLZbWkS6dfqej8g
EsxtMg0cPx7wTW5veSyv+9ONVKVo3d+AwKlryDfPJBBKCh/MpdY6JBig8v5kWllfA/BAlyFHlhAG
nGBBX7FqTD/klvLnb6neg3jaaa2ec5NszDno8VDKJko71ItEd8r9tP0itSOMZKtMiUbbzsR7alne
3InTHNbpferdotjHJQal0VQpiZd5e+njgf976fyTo/xfkk/J9KDd5MHIACK3QGBOhWOjfJ8WyrjG
vGHC75CIxDf5/Xo/KXdQC+bn+XCLqVyfsHZoYDfWdJW2YQL4opyKtNp+GZYU9okVpGm4v/nt9XwS
OBghn3QEZTvwnOdP1p3v52KBqOdmMLWl1oYKYKZYb0HIbbhMGcI2PZ0yeEem8L3/YSpKveHy1tnM
jT5aKoo2I6NeeBkP0qx+InjBEWe/R+HFP8vYmPNC5QlQp++ZsB+Foqp0M5LTSOZ/g+ip09ObOCar
EODeOr2jmTq7U8H600I4N8X62J1tRN3B7m3FQJoaiLyK3nyCe+qQ8DFREcodikfpDNFl8msQg4xm
jWDdTIiqVqPMI894+Ety8CUGbV/tKXLSlKJnCx4zKo2UQqOajkMnnrk74e5HAnMsraNUbnaxKjtk
IZSMupAvvXRPkyTUE9EK56ZSp9JrNjW6++Ed7dF6V61WTmWGLPfefl++jX+fDC3qcvmf0Iv6Z2+n
AiSahhP63pItZqURYJElWw0/Vaa518+G4FvVSwsnoUMlpMDoHMHfqRbQ/BLDFRsz7GZ5AES35ssR
/fid3sOgeWzlS8OLWAb8Ee3ZQoyzxZfwFPq+/r4MInpAq2L+KvGDp/Ch2XRXbCTum6D84fGJbs19
YPaSDNSc7R2eLXzPKekowwDmPsfLZbAMnd2qhf/q7decDIjz1mqGtbIa2Osy3vZtahRz4ONL6Iv5
o7C6RAA403GqABuGDSxT/HUC0cBRGUSB9aZ30DY9mB8Gae2YPoVDK5f853Y3EGiUODM24cnF0Yv+
NDG+WI7ZdISg7RzWYkzqrkS5FmrsUCFhhKnhdwb78lAJmvqfR7ojzAmLd96sv1VWARGwQnXldxr+
kKjd3PtZcs/InNRxYEaADencvWqbS962XPDB092qdQgLuFkZcdTxdZvROiIoAxlqshq3EtA2eBwv
9JsHjxef8aiMi2uh5X9JpUrs/cGWzHJASD8LqEoEPt30ZonVk57AzT8UsCIxBJPOqmadd2I5Y+WB
ak+8RriVnguJD2fJwGzXv0Ko+z4Xl1m1x/e+POCKJXRObfSOjdms+ExGOBWzsO3GRfZtkcr2+zH2
yTP6HZuDYKutOFC+xTVelWkeLpO/rHwN7H8Q7g4PgM3ec/xVb/BofiI74S0o2CJYDu0cS9kilR7f
um7Ou6SCBJQOqoIONrWHEkPQzJQHzI2CUWQXZqWQTAfhUAdNyvzoWBpiifbZ6dVnrcxwBX6IMt0+
tbfLLGVKWE+8ZvNsH6KmSq52CI/bYbCKn008m40QHdNUXRhfGELqPxwoU7/Q18eHricItIXRr76j
ADW6sfJ/hBFCLt9tg2hR6gbg3hDP8xmFuRWIMowFab5Al/cxOLZsO0SqgvAFn3feLGKKhvX3vKQt
Dw7NMj1LaQio4PiG43sIhUpaMh3aIdjhSY6mrFwWUPu+LeY3iQh7uFJ9G/lkG/7jrWkl7G9QOSNE
f7f0xjAkZCVfn+auhVhalnQFFUunaSqBjPnk39MgiB+ort5uh+KEtBhAKWGjcmbZUWKstQzn53e5
k9JFu5Es+gL2IcWm8wWy9+JOuvUvufouoZgSntxj9DKYzBOhjDfw1J53mSI0uqnt+E1+QcGUrUne
xfx4COSSck4zjcc67P/BZTi45v60KqI2I1gGySunmJaVFNlQtXJKDhDczkYq3yAfD5OprfEz7BTu
3+gJJjx6wbnVQ/ab84jJBN3ew/ZGG8Yr2gpy48JEV1/FfaZgAyE+fB4Da1xR6nrlCg2AdHY+29Px
4OkyCGvI/aSIRgW41QG0bQFtpVNiaemkFnwLYCpZU139PcAaB59k+rhI/X67hlXtrgbCzOqe8Ku8
D+72JPq08w6OF9UKSEseoRgg4BRrk8jNquZnlwwtHFdaSVh90DOPVQd+JH/eQAS7QvZoVsAvroE2
eCUoLXt4/aCRUsbbNz4xXvBflQZKv8BJVfZOmQGJf4b4xYlxMaP42ZSZHJ6OqKd7Kl1YGVXUsAex
YB5W0IHc0ROEX4UKf7jCIOgI3XjIzZrqYpC0c86IgpVE/9UIUTx2lhdRYAE5hAh0Ih344fuuPyTu
CEaqo8HQEL1/q3SAxvdvYQCj8fmoo6cWtYA+1glLsS1SjhS/SYUi3zvoUjbGc8pcvzyysD7td6/z
vhCBMSmGekA3zNe8W1KBHjp+m7b9KJIPgt0uudD406UPHIDjFSG4h0m0/jIMBjwD8q7e5USp4d8m
f8gVsfsBF81K70pJWT+vtWTCmNYNsNly2m3cwifTAtu9gvowB+SpFFBQD41TTnK5sdWLSTmDgeqV
Wdc/e/B9inFcckerEYfDh3tRHDITtZxYGn8VN1AtY6UJ/OAIEZSMZe/lApOQK98jfJuLYdFfhrgV
aUDsLZ64FuHZ8UD3BRBgjrcqlae6a+zi/q6j8AI8eMAtB6hDalPshmu9orY9BPvHjDJAq9RZczO4
X/mhX6vwAPoppxdu0NC9pNg1jWYsJmqKegU3a3bCJtaSg9RIZ9U1FxpFcoz8jk2OyHJsMOIzPcXV
HTmslh5HqZLty49bWmCjLKU53fVR2OPuZSiKFqdL8jfbLeH9yTEfH1AN8ZFByk4++yIbAprUmx3A
zagM4gzJRED9tF8Gs1Dz16Z01Jo9UdRl3E/HUkGKBCQG0ZBsvtlnEUp1AX/O62D+6cbjUDH2vdYr
1p028dGIuHhrx1tewyDjutiIRPDcy262FMEdaKEkZrH/aYq8eEqDTMXU7c5gF07ZLfUAk5rzTllH
N6jB4WiEABGt1hgqwL3z1x2xA/o24n+yNq46km5LO8zkV5WHIQ8aFKEWcfocdL4njtim8WDypHx6
tA0AtDS053q7HPbo2ugGUxcWSPoIgPnfksqUi3gbIxFuQ+dB8CUPPGs1aVOzsDUR8omIz9vMbH7L
Wz0s4ZJemDYTXJi6u+xvd9OigJeFc4Rst6ZJQ1LNd8WOeUbbOK9meGMpp0/5FlGtUP1eRc5OuEhi
PeqSOwXGoIV/XwEUZKS3Hp7QfphiW2ZyMFdn0Q58k2AYXN1/HVNccUW3fl4SGVrdTaKt9r4rYDNs
meXHKHFlnohJraZDPO6nxKnVbxeGvElsae9QWZqY0DItznVBSVXPcFeXSYSiwYjH10Fwi8uIbNyG
PysV9hdmpPfqkrcyAiPwJxxb0t5iKIVgjOSc7tATMC7HykR3sHa4xXdJHQvfqKpcj2gF3yBoNPpV
FxWGE30Xx3aURPgVjOzo0fmpyw4YpR++MxQ48vlE77wd8TIir6yhhFwaAdMdbLkg7U3q4BXtO+qG
YcQ8inVnT/6h9SiQEmqp1/iV5LsZTanEfaFEU/hA6+ZqHi9E/v7G9qLoItfGbDupTAfnZVo5iR6r
yi9SIsEZUjxSDRfIT/0M3OfXTwXExhCngiv+uAZLTd5VdYQ45P4kQfkdoHf2zM0oCS3GAtofGXIW
2lkR5PjzAEc6Xz5fy6PQo3u0Ofe/Ma4Iib1myyEcy3d0skyNBHWiquL7sjNR8Z8H/IBZJUQRVt1Z
5aTvzoUYIrr2gvZvCUtcCQcP2oFJbGbEt1COag2FyUqfM+0EyGIjwfpN90cY04pmvCHMM7ivkjRl
s6Sjfs2CIfB2Wc9L6LIi6NNcdkBoR+k1JhPnUTJmXwe36CulK4EnwAABeMzcHoEgz2Df2qA4gbUI
NgnFhcOOnHi941hu7QL5dFu4/SKQWYSYqf6bHidn724QT7eguOkqfAbYhh82+yba+hwHpSp5dscC
xg+hWT+FsTsfcDcKjftzhVK3QCDMTm5nILjtg6Tt7zS/hTJNMjPNrKf9+F/0ACX495fVWJuRNh71
Hh1CiONFPI+S824FYayjEiWvRp9DDUeiNi8GlzcE3BM3HvXjxeP+yFeHkKUAt5VTrBXWyYgb6Cjf
9eHgludtmRwrCLOePgZHFjYzs+LySohdo+ud/rfyQ10zyYNwqNHUysEh8sklTt/o1QhIm5ffZjTi
TW8RN5CR8KDerii02MkLbP+0mQb/qbilzckIVb2pBc6q7auTVt3eTI2VizEiL5l29zkBEbJf4Bsc
ETTN1W2XuEzaJfGOjjzq8/r22DTTPANtUoaJm1dY2nMKPCIuHmAIhYGbD2RwbV0U5BAuwPC6S8Gg
/GsiwGey0CkT6g6NwJPyOwxvUxagVm3LQ0r1HFC4yNClFUwwOJ9v00XIPHGdmcTFqNHVhJpX9t4S
+4JV0OPep5U1QweofXKzDVyIFOsPyatUCMw9utf3Re7Bdkh3b6uPkYN5Zoa8yKMTfhiKpJx2T+I+
NPeTDNul6SYrTHIE7W8y/Qx7lJKPMxJoBx0PJprtkQVWjuv7WCLVgdTFXO1rm1yuIrEcpdN2EYm+
c9R6L4E01L0OaANwNg4q25tljcR8fJOyCfs3K4dyKQyq7I99ZHGJi9PXSXxcv/2cE3W/i+BsS3jg
gDa+pqkw9x+lwT/GPkpSzbIEd21oaHu+h2FPUwPdW1OfC0Xy6oGyilfmGNz2xhyxphx0/B66lr53
QU9Y+oJ/Ua9Vc4yiKNqdSEXUu60NeQD36b1EjDGVTPXvTaK2cWcKwslXGf2ZME0bhSNZzv/sFbZ5
TyruySt1bWg+t8bAz9hClbqEZ5TihStlqayuSZI8+WVEgfoBe38kcDKpSKqOIVzQ/aUNF+c86KnK
8hKjca52pix+vnrngxffJFX/XtR9CkfGjN5sCY5lJ2Wj2Z4p4wCayS9MjCnHEpCvWSPmhpM++ML/
SRKvATyATfXsOozRJNb+0R6Z/1tpcf/T+GYEfRSMD395ATfos9Vi9O+0ZCl5Fxqocb4YrIh29Bdt
WBP3pf6dDqrPhoqE/+gVqGVtvR4m5DTZJmMN+GmvqOqlT5RCLp8+z+q7e2ceTLDVE/YWlap2r5zg
oJplOveVnY3OfHqKhUumeMkINEHRb5IOf88zKWfYZtWTdFie45A1NLqNGKLjIb0Ey72cSdgP+PL4
J3iQhbojT7dmLk+hryS4kxlOd8fxV4O08vVDJpfNBvd+pYRAAsA1pCB6EnwITbKmBw/GHfzRNhtM
d1uaeQvqU/JrgWCWgg805AbAyVy5/vszBBGeYP7y4myRrH75FhdDuUPLDTX/F63vFmhKQfEQs9O4
Y1zU9bnzA4GS7mHqfgnACj857UGsF7pQdv0WQl1WHu2xdszet5yv69HG7FpA/Al/1Z/wb783droG
Dg91g66azMPSheXxUwXMOGM4JLMz+chvyLT0a946Qipx/575WEhlyD1V72UiBNHWQHT9PtO/YZgk
+ElteY6dUbwYydcjdXl4bytYs9KyNi7n5YTz8UzNsJ4Tl/8LRzIlz6OgI5r0Yrn012Xhe4Cx+HQ1
J3Oi0CeiOoOOAADSgznlGx3WbarT/L6MJbtj5zaUGYirQF7XZnP8PjFSrbwSLGuzyKjlczObIA1q
MT6zn1bLrqyNEvNZo2Xp/G+mH86OMaqXZN0W+pJ4Y0kyiRmhEQRL1Ge8Y2zjx2q1H1i60ve5xsxV
+Ay4gte1Thhss3aBmjtG1b84hGa2VGyjLCEYGjSeqhMVY8qC1/ALHT92r1CKLOHE8UsvQXMj4AyY
kgcUssb157fKWF6DXAO71JguwqED8dqC14H4LcbaFN+7nWRL5SldwRSDGld+skVEKswu5+ZewsEK
8HgryVzglDhcb2lnkmJXESWhsctxwpfa+A8xfHU7k1abVgSYWjZ53XkSpdcFam2VUQT3XLZi+159
U3XGxgGJaepYF526/Xz0mmdouosGzruvVIjDRDX1hAXXeskuvw/FF+sHXfITIhZGPmIy93W8nqgO
W7uF/1uHbr6Bc+/HsQdipwCOpJzEbkJwmeEom7JoPSRUrtKMhaJfXf9jFjdxxT0zn4KGHC+N9rWf
jHpQZC1xxRclrY6sjK1CBEcxPsa/kHRbIxlFy3eJhPaISlJ6XOm43qsK2odNaSoVLKzvImiTAgCl
DQMNf912/DaiKgTbD4uPqRBgFflubPY8odoaH7647P6Ur26B53611uQGdSjVmtnx6LLGdFsEIGni
gpDiOnX07AVNo5Mt+QlhRnO0t30iCj6+9DVegAC6hwCFqfAH41KGZFnRjwsqYM9ZVR87sFQl3VAO
o0hnULCHDmIgBM6n9qm3aVgvK+IKDWDv1m6cMAWlFacCUDa6dZm0Te9UW0vqbLPnjF65Lg+61Nh8
pKv1Aj/9YN4i2BHXIiUu2oL7q4vcEKpmScJq3nMkNLvnl0Lsti0UsoWa5Oj/bgKR2+SDWRPnb2NN
l6FDOM5oc1eyj4XyYOATFeShDZDGvAG5eKqFm11o8O4ENy985hT84PSptyQ0e5SrnlOaIua4fLdZ
aoux1zZGn98n8uPD59gElkV1V4AApMRvuxEI/1vnKQE+7C+TJtR6QpSiuL4r1bOdfuOngE20amKv
px0TM/eTX2jLOQdVIjstHwq+nu1/L/o5nf/9Oi0FnXFaIAG1KWIeTSohJGCpuRwxrW8vVIxNtv/i
14R+hnEEvc9ORDe7ojMQR3DrPHPK5Fw9GW9CYhSdclry72CAQBSuRPo6AQUYouxV9c2v54LCHo/c
LGUTfqbnDHA2U0+V22TXpCdyUnMQrDzefcRu4uDebOTF7R/rzJ6OkOgqrvzb5MVtr6VVSR+72M7A
XcNQ2ltzOen5oXErOUFvWEuUwtgIIGlNNaZN2HhPv1dxD/RwIPTzFm2/WUGjdvSfxF5FZMuepgP/
z4z+ECm/CEV5zXujzDdVF7vdBxGVkjQJ3SFwyK7I54U9j2t8lxF3ZSNFmBgSVEkhgI2zb8u7SjgC
VG6JGL9AgwgNP/sIceHkURG/IN/OvBlCxsuGkaS+K/5h8izoZ5/l+E5CzcIrmjF+wvis3VczxkKR
BvoXYOGLBumJS5UUZTw9MsyGrN5FHoBrKdDF2ey+6MTB11j0wSYHxXONqBmSfsZYXw0aAEfjTFv6
0+bcE7kD6VwmePrPK6OrHNodKtW65FWYftg/pSHguwsi4tLRp9Hr/agHjJ71zxyYrAQj5sCFeAHP
JfWIW9jUIWBxOrcddBNBgi9duHI/uuWmbYmgXIFmiguA7ocxmO8R3/SaiDkALtinfyaqZYECYh5T
ERMUw/rwpms95Em4D9tT5Jxb36pTcSPyvNlXarJUKPIf8Zb8KF2/2cDQ/rpqcRmEWsQFDkImXlMZ
MR3OMrDyXo6lx9EN5BC6qtRPf6JQS6C/0QT31eio3oiQP+1mXuJ7vMGOfq+rSAsE4NOEkCph4wd/
CgAXWvLAi7DgXP0mMLyejKxVEaQozwtdJQ9/rGZeOuU8R6s233qcHmUgiKeSEg7NVik52kdQb77B
JVaQVfS6vHMauaVlMNDvIoj5jYWWYm/iwigpwl9QU0HUaGpjuTlCzrP9T4NE/felkaT2XBj0OT+I
oQNoYzUdTc6s6LFifm+V57XUuzUkcx7I+RG5bvQ+vMUlcBXwEjkxjrFdMps5fyYG1oatw/SrsGzk
1JRiYXZ6qQTas/+k+HE0Ek0FRcd5MCzdnbeV5iRNLaNQ7YsCaSn7wBlMarpFSQ935OIv0AddpRVh
+yE6b05k+Dew3jt1c7j/CNwI6MvRIvUuR31YxdF/p11tZRt6GN019Adhw3X908uFdvooDziB4F0u
vD5idVrziqK6hf1gMpcpN1YKjrWuNI80bWKc9i04NPZX/8IgifsfXfrJ+3Agdt2DRfUlFMjbYwYT
9sLCkxSgY+b8pSE1wuGPwbGiOWiDY77sYbQXUJENbsGuMlZkRe6SFDY3EMgYqGEbMdqfvHWNzvjC
nTOBdCrDC/E7r+cALC8QNYfkwSKHi7iYI8SQUJdTfZVJmKVios8c8nZM6c21T1CKQqh3tSQZRvUU
HY+2dU80afSFes+gPi+2miXwOPpH2XGh1bkZC2IT4T4D30H5jdfSf+dbw+43CoGGvnE19ZLDb5pw
OB3jZWIvrMSDJB8yT4EH6Tu2L6U2kipc4xz1F/SEmrmNPQpDXBwoQ2OFd+X6iySVit12kOVb0mWV
gW5kDCHQ5f0hC4XOhqj+Cmfr3Poa9NyFGpy6b27XfuYhI/+YAWjaJrO6F7Wue5IJCtFwwE7CNxY2
CDJb8mIvhxCjSW/r0PbElTChtjrUD2bGEANBmENC0S+aKp5p3Fyqx2HuG+RhsPiZI734sprY12mY
guWDAGttQvihOglEQWirXUtnZEvaJ1zdqibNq0ZZXMTBv6GUvFAQMJoP0BLpx77wEOxMJctXjpap
S/0MtUoK1fSzszIOUn0eO1lNgoDpBZ4U/DKdt0eTacH3ZxqjDXrLdDqe55Bthog2wLpdTZ5AuUbk
LQZny16iLh2dfgGaaZ+6fzJwIYLNJJTTwMaapVqsUHnQKDIv9QHmDWTXtpTV0HsIBcT0cdoEH4hj
+RB7NpuxsVhubCbSZBoyqwPVA9VTvD1yH4Q6mQWiG4vpfSkfM4bAg7WJ0JihzFH2S/tc5WMCgb0q
D56zHZKiVIg4JxKO+MqcZAepKF3wPPGTikq4Wjj12PnP7rrfONxklnZ0fS3eN7Sg0ARTVcBHllNF
8bA/u/gvw86sknNG5+7ZNPzzf3mOHvgUnI0NikCgjjnidRZ8kkCuX/NWzzIJHT5w2wzZ7IYplTF6
Lf1KnPYxeVXgvW+ItKh9eSW+wW+ZUiGgeqhIttqu71GaNpXqyNgjKHQV4KsLEEIPh1KIQZkjq35h
ZaGD8oMt5qDEKimF/1bfsttkzzsk3Nf86pRPc+TkF09alEXV3wltZCgYmhdwhrhkUrXtxwDxA9Mh
VOmCHyhCQwA3PbaZIrGPsRQeqT4WGnJAh1bon7VW2jbj6+jLuzZF340Jndp6fA/0uiui5x8yDGeT
BApGz+KVhky8OS9l6gsaTYP3eaZX9A9DbqYtuCM/r5N9K/CPy+65XOZZf9fBHBEHqYhLsfinFbOY
GwVnEQptx8U7Zco74iw/hv5h2c4ov76kF+gmaMK/N9YR6W47UXQAel9uY0XJBdusPRMiGRFfE1qd
r34VLejI99q7wOst9l098JpV4WEpQTqC3ig6vrHanfP6+0o5KVGg/9qZaLRixTTef1Bdv9Iyfkoe
DOpWt8X3CU5vCwnGrUMfniFfz6aoet3AbEfCyXKvkKJyuhODEw6RlBppe4HKeo+8lReXLkLlx8ZB
ieBDLnni+s3De3Dcr2hheAkyjJyEbHWw6KuYjGE4cJcX4BG3awEvLDJX1ScliEC5JYusf653YdfH
ct7Xtf0GdPSTl37+BzUPsfW39/59ZV5bD2wywK7VykCcVcBQJvh6IYdj62W7IKl5VAx3OcVy6M5D
NruAPOi5ZkWZypmS4S8HBjHuSVd1fWb6cc6gBU/E2xg5aWGjJd6Nlxvdki15KY3ydNEqpN9x5WPG
KvaIEzxB4Xb8qgaH2W7WEYXtIsOhHLQHgzBXl4Nwqe1Tqsua6EM98HTT4ilLoxl1TzCFX1jVGtER
jJFVZSvomML8r8Ag8ieUg3WOScZlwLJt1Lojj+p5OuX1tT2CA4UURvIOT3LySTsBzFReVfhnH95H
Z7g0tJB1vtmmAjUqJiWTT2DoIWOatJiboeMTqioZN2zSxKcezzAR6XF330QqJxACx/F8xBYfzB7C
83r/jHJsa8FpK86y2c13B80jbD3JHCnqPtvDmqG7IZQNcdfVLgf89yA3sW3WjEf0EQn/RPcODCKg
eo7Mv9QwQT1pB63T6nrs519WfgGS4UfoO2sr8PgUzbYTsmamODe5Qxr1ZnTdnNh63gVEalL/FMjV
44bV8qZVt+pqqu6HhPcaH82EdSOqlXAO3ODCmL3kQ9HDu3h7O5EevJZn52amJusGMW6J7OuELvZ+
+9IdUIrKjOBJGl8GXEaIevX34o3ZaP4jVGc+iXXCjTF9viLR3XpZH8uhEoLfnzMY7hfU0yT0rIis
A5lJjVL73+XgUqldeCkH1JTrNXAADdCCqoWx33cEBsIs6V9AnjWIJ8qi2XOLJFyAkUIhmkyTRjME
+TZZk3LtqKZdS3D2EC7RZbRjAcWn2ObI+fqntD+Z984qQYFHpFA1aXbO6IDBNeozxxxiQ229ucEL
SGZOnzkdeCGEp/rodkQcUFGUZ416VrrviBT98X0chSCX/c8VtdxwMTI1WakA6LXs3094Mum86+bC
OvqzgFrMlpjYdG4O/lqmP8GLNZ4iL8P1YwluAt9KhqpXGLg4GbHAqJIFo3fxicEsmha0oUd+MZkj
7Luuyi+Iw7A4u0GqGFfIqG5brQbHpKbpalLg3MhsUCnm5hvEXb/OkmAY7aGykjt1AyhF9QHWmUQN
Oh7xhfSxqXZNdzFLhYIbxPtCQ/CjKzHvfNzWwfpW7eKQunrUxk5x0KPwhvwfsvV3Xoj3tdGGdz3k
QUa4VyyOzebCmUFIEwdoqhn+pBHCWd1uXidqoJSY6+rsYiJe7uvCwA2RrPwDJ7/J3gYGEU07vOOy
JB6BBTArkfcDYx7FOsrW5zbaq+fMTa1alXxMuXwruX4U+uxVcwt92kTITOpejs61LFwTv7CncO5+
YfOF5Qe13wb8X8/VPKukzlyqiNzF2jAKS4LjxBKcm5fM+k2auuvWT2ieSRD6eJw2z+tnCelE172/
MjTmFhR+11epEW+moI89vmi4dZ2uk1xFzw/vSumFlta2K9OM5DhqNYai9efmdHmNGvq1Mbc0m5N6
iLHXV9LFHqGtyctouBqKyo8s4lgny0KuTXBxTF+V9Fjxuh48ESrChHhQSEtZ5/ooeSYKcFjyBdqw
ffCEBUA1that7i79Aj+b9U2+4HFrSGVIklUahtb/7sMJaT9N7eNomDWHnOHVG2mUPkmTGqOIRdEo
182FTdM3x0J5j1iw9ZOE44bK6NXJ6jn7gOdtTrExwVNjwrAV+hIdjEz4aw2bX2RKiAiLPuwr2ygY
pulcrJ7xQloWwn40zwqP3SZN1kVwRdnW+PAsCExZMuOc0nnrF+Ius0ssHohckGqK1EJDH6YHuGRZ
UXgC6QsmnJVt6Twx8YfOuQ/Ke+YJ1N0tj8XHj1eQY/4C1Wo4nORJkvcYLRCR++xHT9DdVl+/6hOp
ZDWA4TSjl25ISPg4UWX/2vrayD6ajMZ/ezT3pcUzJ3GmwhnsvqiCH2ZT4q6FzLSVswg7Y9fDi+9v
6rGoWZkSAt/WqAKLjD6TEQsb5Z7J4BVYbJZc9/amDFn9jMD4wkHm4b2NnpGOedgY2hqVpltyJhM2
dGRgjF4JOoCccPnWdvg6QgZ/k6hcRONEDtZrYkkG5z8RLtmmu0ZyN7l5Zd6nk5+r41z3KcdS9YHT
6vl7mkHaAAtI1L4JdoXPNFaZe5nlDNKHipLbIKVLFrwlhZGk74e2KIQ4mDWZO4vljioKRQf375jH
4LdqqCCgSmuZaQtZfDFqorHZI3DhC4mLoCoc0SdmdVHUKcoLd6U6Fx8vjqxR7WdvZajUxMAaRgMV
GXQdzbHHGDdXw7n5V2KSO0Bep+qTRmXG/nxVEWx0vger5QB3QLzqb9S1nZANNqh3PWbVjK3Byyhk
aYHKW4b/yfBpmN2YLvhcpeTb5daQHIu5qfqzcmfEJe/Cw9YF7QfiGYf0z/hzcy6vG4LPIp8GXU0F
G2nBNyq6DicIWLt3keiFBcTTV9EIswXZdXryc6nfuVu3xWMz7t3zuNhtK/G4oGVJTq8hUDTUFC7F
3SEfhVgZ0/mkidPUEIASkCTYE9f/Z2PiN0fBEciwy189QZR2L6m3egqIbV0rmWk8+Q1AfBkJFSwp
kOX2tOKXpix/J7bGqxedkCFTtvX0VIOnaZ0yeKjeYf/fudJxRxokV15kOHhUnPTaUuZzeKw17J3C
0NqdcFgsR+ePuMY1DyNfosRTIoXquSoAyo2epaoAGNZFWoIw8N9mRkGH1euOk4vmD4BtM64BPpzF
7XaHb9YUN0Wb/2s7RlGY+UUtO5Pw05hXafw96/BxXyE9wSEpREbv8ffhxrR2fGE40e3HJBS82HZr
iQdOmXJmSRV/2f/Isbm5v+peWRv5sGWW8Huz4h1Q4yLz5EEpuwk3qHkitaevqZZo555B2xvXftoj
op1Wv64L4908PpKXR0HG/HcjHKdcCU7ckksVEVqRO/g2XXyFZ1hvotJZfaz1cSem9BlKTfPRXvnP
4gkYgye+zeiTD2rbRVQGaCtGQcF+rVDY1tzuDhIdXWS30CgH05EKdj/rWtlyw/YOL69XFdp15a+O
y3q3LjfxMQ93f65zHyudk8wiu5J4L0A96j5xVFoCG3iM+PM+4hN+q69e43WsYUMSKvSeyNDvfr/c
hKyCr6SRl3TVSqqBWO3WhBpcxT1WOPr+sgt/b9v/QxXZajAEdowz8DIgSIEITDbD1yo8p77/2Bya
242YmOKaQmPyxcQUTaGeAb02ghli9SVM7e1fFrmPYkXz+Aci9zYgrXhIqpVdwZPPUTH+wOq6i7B+
o3KK3yJ83b9d/kYgfXfgECUAs8afChCB9fnRHJLIlHlu7mNgJeVYBjmySrc/ipFwtvlqYXoJq238
tUP4tmOpnGjCMdnMOfxAm6R5LL/GhyEqk8XZnMgRNaJlCOtISQfGpkr4WUVpMy20qrM8yLABP/iw
JWo4DpLHZErxZrV3ft2Bq+o/9tmL7CtxkA6sRkLsJ/SHZ37hORioZpCuWhvVCPookQkCryYGmMKH
SIkOBzXskpnaZe9rlCGt1jd3dj+7IVTJ2RX21nNOf+NZSMejpY0GVdxOT66+z9sRzBkDoncnjbfB
b/VJh3VrES6qm2cUaV/4SvzdPcyCMnVqpuitCUNO7dxvqKGVbemfA6LA+iZ8e7HmfDsKEH4Zt5mK
hncPlX+Evca0F0aeQec8UJYxJ6VHkLepiY4Uicmf1nrq+FepNCm25IVN9Qcc64J2O1JGCbfM+CGv
sQYQsDMlIgp/KDVAVUIemX9MMIp+YnG3g9vk4QE1kw8IeRZJdSRgYuB3CxY3T1zgdD6Os5hHcBcf
mwvrS49RV7thqOgdVeMldnyPhLmkaQFgWyqoRTWlOP9IFC2aFte7CtD/GDcwLuQfFeGMS+NQ0qTh
G1lam5ItCY1PYYdGQRj7yqsEmhyLPGXt9pG2XCtFcJ8fe0NsM5873rSNHROeh9JkrngrQZtqzE/W
AqWfkhgnOM+8FMcZm+tasEhrZY5yeRcYoTACH6jt89OwqXPj7p5qEbgPSMhmJ7JoEHPgfU7lLG1w
qrI+HtzsofdFOTQwWS5MTMni/n5+2RNO+7GSaPROXkM8gbGBMOV/CNf4MwwnFVIj9epzsn5ZHN/C
AloFfOBbZXqboxs0Ae300rt05yTl3ocjmahQvEn+03M3QRlkM/65X/pXRdoimTw6eyLggKAom7zJ
VzRxaCpdkHGCOnJxxcCBVZ4/OkGFSwlwemsvbGh2xaPOk9weokzjp+gIQYTwLGzc39+CB0ewcp0Z
P4BnFYFmOs8tahR3x2bQM0UIz2Ya0zTN7B+vATA2YiqIgwsVLFFLTbWZUJZk558wlasOMzzfcoAm
4Smq6PHK37KJ7Gbp/I3dXnxmPlnqbv/uJbquv5oxOc44jvIJ6nhkEJdUIU/IRnn0LEmmmeUg5WxC
LN9yhPshU1m6s00gGMiYezcoq5NFz1fjQTqG9UXGFN72mQBKx9TAcB/oTjN00nBdFfSjodFvGeuB
HhC92d8MUcoGPf06MGjPzxroIK0kn6J5lOolbwOYjIPRNnhdBF1504/bEj2meSoPCs96VMgwLBEJ
kcRjS/iSQcqPadlZl1Qc9D1d9SGfxgKiVdaTzcw0/vqhZ4r08GvEGL9NCaYZPymFAiLmA2Uzb2Oj
1VadpL+uacw7mqrIaMXo9U6hUAPb0TjAuII7jbseiB7MDl4yCvTL1pyMCxjFSMtInaPnSr/yEbR7
9m8L+7HTgy5eE7rZe4hR+lQ1n8Hn1ZOdGIQx9MqnZNviyhfZiYQnpxXRwW70cGkBsdJ1IHA7IIRW
bBaiuBLUEdhLB9tq0ANmoeXMzu+dYwYbR4XRls19kj8KXuHAz2DtLagfDmJUWbzEbS0uRIiw3M7h
oVhIWudxttWp3zrOIvVoDEX+t+6j404jcJDOAf9C80Qe6jQ7BYwncVOsJSqV0ITZnSZOwh6KOyPD
qmyMygCnSRkaowwdYeFvXdL784kAJUjJIgHD9o5s9EkveOjY4+IhyuZBcenB7OnYhG3ENUBtstNy
0+Z4i8VPknL4wqjceoJLHW9EKjIm3Ivomun6UW9sa8Ol3mvXxH5x8CDjccSk6qrPh11xy0Kp1XkZ
9KQuOc9SHay9qgsU7oxerIO3utT9+hdAGSshJTYIh56JGgFfaYGIC1JbEYPq+KI4a1GjL393neZ/
uUQe5eY3Drek4qDrNrGdG2fb8F1R3mljKG6QnNboSsrv8V0Cf8gQZ0Qqxj4xBm9V9SmGm6tmbcI6
f9H6sEaPK3A8ABnu8qzWErYmzKpjiFq5eJayf3ftIuAiDiHqIZ++k1d4VzpAGgaSG54GuvjuKB/w
JTQzb5QGeSC4nzV2Nq/6z+Tckpl71HSWt2eaBoAUF5klnhmJ3VmqpcQagaYwblcY94tLHBAO+Eeg
z1MzcnnmKqkG366B+csZxdfkfqJOCpvcIzKLHyIygFucwipFqXbQzL1BkZApifxtmTKOyo/JVZhO
x4nQqs+3P9NANc6Q3H+w7ltNX0aoKnT75cs8xVO4z2pQXhFj+4jE3y1U3dnu3krSK5pYnNdHsQCJ
SDypvnBaLKwQA12Q9mA7ZFMBB6DaNTX7zKvRt/9QqL5DvzTmjYwlrgVf+rjvNRjOXh5aMksqshcf
bp/tuAR4OAhEk7lrhnOk7xQ57GLCSusIy7IeIfoDC3hFG3cLq8my3cQxm/tnmK9xc6L7d/q0DdjP
9VLaQj2ixMQV/xYhJDxgfSwr5tURxpdX8quF3L+nd2kXIeHRZEB+PkNwgmCsFMHBHSPouiruE6Zq
JxPY1nELQ81X1rmKBs4uks1PRX07Xmka8W2SKK931xCfEDcYFZt8XyNodOLAbvJUohWrI1L+rTh1
RpWEHcfLnShSnlNNderZdS/6xmniMRqWzi7oCz5KBr3czLZNSb8Cv/XIU7NdTKoE32qI484xVcUx
OZ/50tXxiuMLk50gv1H6F2s0R8ZOqU8P1NghE3XNAPgNG3YTX4+6BM3yWPqXpL3rE0Sf7cWwajs3
fSRVzGRgNT8jT1J3XEwqPBY/NZrzNJOk2A7mvkMmMMzKrIvebE6z3ucclWVtpPZSHl+pZ3/Juv3C
g85B7LfuaQ22pvROWNFIkff7+KquAT+CebJ+enVAGgLw0koON4f1J/RLO7ILur0U6eFf9yOU6dzR
HJQ3aZvM33BYwWQOpfV85ON2rb9lfazXQXmnnsALxrtp7PuO3A9eoOE18hD1jJ+nWmtM04fi8f8n
4cDhKYqcW0BT7+4E4T0bng3L5DEcjXTj/qszASiLd7lq574c/uUlYRWcfbu1jEELbagh+sAJCqem
CGBEyzFLArTpwnWQ7BAnl/NvCtfz2jMRupbStZzqUna0JAumg5llC+K9bp2Bf2qMSnnDbruUVz4E
tUQx1Z9kfDmcunN1kHTKQnVjMSNnnhYN1GLx+xZ6xlzdDFXE6j5I3rWN10lcJzIbuXH7wwF8G0IL
hKEukP8m1y3toA14+S4R8aopxd9WBW4mMj44YazPcCZMYoTujWqqKojEJpMapiYWl24nBzeW7MQg
apPvGfkJ8QopcAex2YaKLuMtwVviY6fsY3oJVu/p+hDjS+jUx0qj55zlewYroHw56WDrzA79iy0G
X2dddn0KmhQ2042h5FEG5icR9+sB3b+X6GE2VFgQ1RX58ouaRkMwmkuwvo2vKny0koM60irqz63L
iZbwMQJPLlDsxmclp7ql0Lcb2xIArPK8L3jtJmUzQd3Q+DwMB50EZG8L4qVRIuQNOkz7ZieVYDLY
tFhryzYV3l6zq/qajxOi1JDRXnGCNsPx5J6D4bj4K7UYnW/OZZHURL8O0oXC9SLCD44gJXUJ35aD
TRdlyUQvFcGyaYHD/0nl4oJmVbpAR1QgjyI6POigTP2fi1QerVc6sxvRKZonE0iTIio17TV9s7CT
i6e9DOuA4SROwyvfjqxBhd9THNYkvAlUSN0pN1MpH6pQhWJCaUVQf5xdB5g2X5O+Rl4PiWpj9J0R
rRKdTMOBqtgukJYrOeNQujfVZUR0Q0g1mwaww+5Za2XtQiPQEBb7D4UUzGulyJRV/iWNnPTBFgeH
JsC2yrDqDc+6Oq/9IiqVer0xFsVX7aitbtfvTG7PatiW9To1tn3jEEPvj9Vu5l9A8SCGGyFxL8Vw
EYyPOhpk0fzrhFXI/AyyV1scDgL2iFby1m6JALC0FuZEihaUUa+7i8MFKij3nKhqndoukwqUT/VW
UmbBgOVnT7ZjJ6d0qWpVlM9N3FcfZ9sLcjKpRWF40WYXhL8DPa/dPhahyTi1kno94sOVAZjvprku
35I2I2J/MEeGPHTup2rPA1mpaCyzcQ6A7yjzbI7QyQIqZeFmgX5IwV2YxS5k+EM/6/n72jQj5h5R
B4LIJLz/DvW0LTpQBHezC3A2bRvDyUSDM9NXfthCVIbog37Oxyy1RwVbH9oJKB65+d/dRZ4JJv4k
wpesrn3xHjlQZLCktuIjNJmcnaxze9Hvio73+yFeEbB7RvR9tQfrSf1rXkGtKp1X+ZnWCQ2kqqzr
EVJxXDzUULtllrHZO0CZdR6k+L0ROAILC/2TywJdr0v3i2+lZ0nz1bAST3z5RhPnFHVL/lQtFJ03
MwOCYbDR7PGrAESU3Z/PA8A9qEOCCKaB/jbbgbeNTtDaWeJSAYKDgV8rc7ogtsnfg976QPZKg/8Q
534uohCVMfzC6ZGbFjvAni9x+GqY2L/RYTYrBK2kZTo2wxdF1JC8iDTQaUw2AcdicG44WDS02N3j
tBZOGDx3oUOL4HAsxtnFD7TfRR0WvCJooFiIWkEStCV8mL1PjLwkTOm5KBwlcNTnx+SO05kISxN5
cIKGNkMXFGRj3FzzQWInEan7SEs5pEHcY0EYIeb1U7Qsa6omvZJCvkxXem3YHBsrLZbYbLGiuSUs
6Wb+HsiYVgujZFdJXVDV86VodKtwTfV2U0Rqyc6bQgt09qcmOQtqvva3Oib8LJB7gQ25tk1XmV7p
7ciQh5FRKzbQ0Vz9p8u19JmHfyNZk6CkUrs0Jr9N3A7d5ud5sjFYFOcoOYXiu9MhA+MQNRBlheKx
VEBKncxxhWJK1YIQ6dS8v5iafI3IsHtpokHZhYw0ZkS0V/V66AxXAVgsOOA+NStiQBlySiUVtvx9
/vpFQnx9i0Bh9SK1gNC/5rU62A0S9ARTo32GR2cn8ny1+11RTAvMc2GotNSnFMzpxNMTTAt9LcbZ
MYB/RwhVBOzhGDBr07amlwCmNyCVM2tECHBpC/7PAwc+V3jpejSlU/5UAurRjII3lZPLwhOlOt9T
YTM2ykpekzRKySz/bSI5nqjKZ9MBNKKdm/q6be2SPt8/Rs7vpcHb3kjrcYqDUFBzRHOAjMm1xFDg
/roBWT9mg9zF4tN1CDKT4WwKwUyeL1hduVXoNjtAYceZr7b90ha9VYHb3XmhQ5UItvApmkX7XKMf
t0Han1+lIyKL07qFV+/duJCIIbDt0i947k9FNc+oHR6/KwqJI6QERbtsY3Y8Ni0/j2TIpkSN4rhY
sAi9WjEpKGuBC6e2am/BAoMczC/FnyUlv/JpEeKXBtqRk4k1TkFnjLbKkIhvEM9+k8AVMy+Mgqah
blQo2Ur2tC+TPj/8XH11Dli9QyRb5T+MKrDqMFxnQrpoTgJ0caGyMptpHC93pES4d0Z+OLDiV0iB
tcFobw3dvhVhefHtSh33wDFy2nZ3mSYoHCwLmFHyV4zBXR8beMcf+neTIlcqmuLVcKYrzaynGvVd
vtl1XH2rIM6UkgmEfnKtIErYqEPE3R0GcqjGDvM4j4T77YjLVl7QSn9EfKzA18V2NeCdnkVRHArj
yqT9COQP5aQ62wmDwCAY16agY55X9Jz1WGko9VNpcTrvFmQn4qblcN5Fwh/GjkNZrFACF4N4hNrg
3pCvKIKcw43mRucKkS7rxQ8hCuIWm4ZZMUzKGTXazX/GTXqqwWItM3TuchNtRZtTQXUluOknoHb+
l7qtrhF6ZpDX9TMiMHk78vEACDegCApNO2OJY+vtW9+3MIsdiZXv6mLE+YlY6pD0MPaR1aEy4mh3
L9o3OfgKePe84TL1qFB4FT6+jntnlVoLYzKVMsXDiWZuDAQlZFvrSyHJX+U8HmQz6YH01rl9CbGo
0rb+VL2lWc2v0/yuFj19uubbev27p5nFLcelymdyS1qMvhHfSq2um/vNbCDcUPKf7P30bDjLJ0sJ
BXfWq03Rc9/JC6TczRH0d3tGMayJdYE5m8fYKPS/ftfDffVTiagM/MkGYQM5K/CYc9C6kfZic7kh
L3/hzBBJw3fLFngSWTQxJgVF3W58LqI7xGIZfseavuGYILDVsZo34wFFdbp1Ty0UsGTsPkwPAIar
zQ0+LDC+LZ2SnYVq35hBnnGDIW3bFk/KoYtgeo+yA/+vXo+PEznBWNr9XIzYcK9hDFqqcURLBBq3
VpQwymCa1Pdd8UY1FU6jfVH9v71CmOfOM91UtMeGuajOJgMSOkJnb4peJytUXgeJfWyRdItSfIry
NpgGBoib40lmxG+TizemQmbTYnC3ID3XRP8Fa8fcpPJhsGtTSCqwP0Sm/Dktx1W8wia0jkLU+H2r
CDrV7NELxPahhP4xuX9uURcMK4t8Zsxzq3aw2tQOZdmfzrj7mw2pqqjXtPdqZdPdtBiXSzC6kj6E
6b+0+CyqJtw1odO1k+UnY5hzC6/CJBRDfSnH+Ya/8YvTME+ori3oAcKTpUAFaYVgP5Yl0NQbQ8Iq
eX7GVqhq1tSa6NGDR71+aPgwfo3RAuYxt2JNv7qQEsthyIe63FxwFBegZIicedX0QPHxYj0g5NPD
AaxGwhwLHZi/7fUMH64TnjdksaqNn1gN32NViytndmNjlx8fSUpDf75ZiIpCAgY/7BmvML08797S
mHo6Y9OqO6iXJs44K8I+EDoO9PQGNPq8mCjvt06mMbpdL6S7EMQQsd8bshvnGQbFxVTVjp9lO3e9
Nomh3FYK+YZ0p3F8clP7HTEofMGCviBACqTZ9QYponaJo0DxNqiUSUIRy0v+1DAHooJtUuuXE1XH
vtzDnNFpi6DzwWMgTCjipil6H+wDp0IS3Qp1HbcuW+1Ch1ZgqbAgqWixWX/1Mc6fqhuk2NnTtTRs
o184/q760pb1uM8hneXquWLI8Rc/UfRih7+VJes9OihBRSbU8xMD7FcSKZLatbZew3AjPKXwE8Il
iwq+6AtC6JuQpyIQUAf/XXyyD+NLYeXCZvEyzUAgMLeoVnFgsVFaM8b3IS2ykHSM9jltpWU/tXC8
9BPRyb+6YQ6rPGSIiUzgAoqpx+gLzhYtK3XK52Jfrj5eWOHRXgJhvIHd+Q4ikJShdmiX7ahEo7gl
nSgCwU67emleZHg6q/EHGFDAG1JAKQsTxlzvC7YaMesJ5cDXkq6Jy9QUK7AqDO1xm9Y20TkswTqb
M9ERsCS3GnDLahnMchw6baZaspdvt4gKTq1u0NaHVjHEzLEEwJIXSUfxJTX+ZF0ZZJmQ0nyjjNuv
gsaDg3IubTZDAsa9f8QgWQoFhu3J8h8IpwYIK3VkrtNcRb0YIcinOoE+aljKUaWnXWa+ynjfTU4T
TAbf3VMNdpmM2U/aY6wyLJ8ILsqydHc1y3bfm1UKF75RIgENiRmA/yfVkqxCEwJYbwMb/ZZY9Ahl
VXJ7A70LbuKXeD7yzj5sogbyZFd+yG9MarWuK+8WJdA81qTgmyYvTRTzKhVz4xto/7FngDCfhXpH
3m4Fl+V9zF0jwkAB//yYOM0D7qAXQwnnYbidFDOd8JZ0KX7TyqEJqhXHD6TzKSPHQ7k8z3OIMTth
mIXJHADtiN6er+kI4JdulxB7PU1uRoITOU6lHyKinxn57bktuOF2ycpQftBdmuJ8D2uV1kxnC+f4
Cf5WecizQRQXamoc1yCio3eQ8BIISCeg2x8zeRmWmzy2gaRuBxzNfSI3lzgBaYxAtNdjX4mrBnfh
BeEhNZJJLM0oZnO83PN8rCKpbcxa+Xye3LTS8dAXl0ImMZC/eRSvnVV4VD5kjANcBffkVVnQO8C1
SZfTLRYnva2h3cG8RaVz+5bBOnY2jNm3YIqklq9iiP+CzvdlwStqnnvl+sSB452+Ta+GS/M0tKBs
MbDpBVJIHJltOX5bItE16eHUuow8zO/lOkslWzXxYrqa1JDQz12qh/UuouEt/+6JHueK/KRtOtRu
zSXBxiEmQGI1QRmTyR4ICnvmcpF7k7F72IC+HJfahNpopsMBERGuC9c4NYpoQ8b28eXjV2w481IB
Wf6W1EeQmvKriodnv/vyn0sL6H3uAn9Iy+Z6KOg2BEY+/44oe0bze8dDj5dYYec4TvAJFfomLy5U
CRxMwoByHVQI4Su8gskagxHGD2jLkq0+d9rmECQwZ71ib4CCvS0DLv7/az6D8xF3Yu1Vn65zitEn
meRSJ+TI7ERKGzPdStRsBNfblc+mym6VxO6eTUSCtgIZAA/4KMPnAhwnSDWFa6S/zfunwhPo8NWX
lA1/rz9jOwei/CiLiKxUy8mIsKcip6Jjjywl++cNTpPbSOFKXZP3MwETIu8Oc5tj1Rm/HlxOp6ES
7s1V0nndEs2S1TgWqV52e2r7ySTk8Zv6wsRWuI5UjGpx+KYXZx/bx/HbiGAZb7vHT61CYeLVakK8
17A/YnsmYwrvCl69+1wrrHzcQzgzlvCBKuf6XNcrSzDSD99N/PfoNREE4X5rY8eB9+zoxwfvpgR0
u29KOb8gTA+JrYxOsK+FrM4fo7xTkxjX9OejslCiffYt4SZ621clu26LwGNBOmVD3qeRUHPWBhSg
L4I5s/HimzlYjB7awaAQSc42MGP2dzVaAdzuBhU75Aq2/ZPdJje6EIS6zYrdBCMxMqrM07eO2G03
gibqb595taucL+cZr5/A0o+vpvNXipGcMRO26roW5KIupClkqD2B8mlwgT5jV2ljKn+pi/4pFz/G
ruenqQNK3B+1DrGmTikXZCgJBqhAyU1I2Uq4nj1O3HUmlLterZUvFEpFztbhxvNfAMlBtnwDAtvq
+HDoTID+OTfcSVBYDyqcygXfgcjS9S/RAXbCAt0QA1kTo1jnHcuL
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
xI5rRsZ8D/mWscsXgMgqvONi1IR+WUmvlhOeHpoqbkmGbmmCKddy2Qan/TbchxUow2f4O04cfAEu
JYQ5L/DafoWEAHShGyHztGxj4EyJX7x8yqtcAWwgcJlMfy/2Z+sYHVx4ASnUNZeQ8HXpWibYIZuP
FjkTNuAr1SrdQnqwhH5cviaA/5OheQSigRQCP8RRQlRyBxc+biSsCZMpGISZFX2CZjSyU+7V2yWW
ay7r6zDWmMmDZjudTCI4MmCNXIWpp/bhBBuYrBSF+L/5EsYX/jb3bbE7tKSBxKDVS/NsrCqqNgPq
LE6lSb2eW+8BDcfgsBxnkhOXEUv0U/y1UADlGQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
kt+7rNkOSYrcXqbgq36Tjy1mVNbqyEaJJcQomY0hj5jTsV2loT+ykCqTokaSF04RFimKeTBrbOMs
fGmY0J0Y3FLdb9mRm02LfOxlSlD1IAUzPqmK1XSR8d/4MtempkKY0sPLjad2NV3YwFQOuIgbOEwQ
WJexgoWi794m/yDoUFziRVt8L8gAHObe8TsXdCCkIFw1w5BV4qiVphOfsBcAFfGjk1h0eqKL4hHd
+knMywKT44w7gE4DaneMKpcCfQ4X0hNR6jP67PdO/EqqXFjgnAn0wypmmiFT+lBYDb/eP0n/hSzE
W8aox1YjaQtyA9zwXG2XZMpfhHFKcSJlD/u2/Q==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=157728)
`pragma protect data_block
MtdCuyRVwVMltNed0W9s963IEM1TOevhHDGLBM1VnDmAsPLBepDiKwExnBgdfTX+4mBHLfj2CtLh
UNTEX91wFd3OPgNOeTedydghDsO0yck8CYBwzEbc5mDW1HOZ6m2GFR6g1hXZTV4tC5pzN1dv7DGc
fyg/o4QCBi8Rs+CpVC8mLW5mVQ3JryfoIlU5PvdlgQZpyCzVz/l8caCeoPnPkbpVNaRm842kWmgI
sQ7kXDsKr2XHozm7y9YoXy4waUBUb/0XM/fo4map31+pv4Af24tjUDprGbowx9s0ck0cidGfq0tF
mLj/lefGQhISo4WHCzpORN+zRh2RrIiwohTwXu/Ye4fxkrXBX5x9wxhWTIV2Pnn21XO4SaQq65/W
/rq+W4amKjPrCvRLj1VNseMiExp80wAtLvokmVc0LT5gFAqJETfF1/UE0+eK1NrGC+v6+RXQJGaF
1wvXw8IH3F4KuULbnbnX0oD4MwPbkcUq41vxTHmhfM54805oVsHSESMa67+fiLhn1bVx/eFobVzU
1eA7etG0i1+vrFnj8uBCoK2Blfu1z8gT2pGKT05eqoitXi+hiOcAt5+7zVXJ1Cvxs6Ji8T+1ffRe
EEbWlsdN0OG3p10VSH/Qm0O72lxf8LCSWH3FQs94onWSRSjRKn47oWBJ6xw2bcyJD4nQOq9Wfa7F
RI2X5lT+G79547gplCtWJIQPagruyWwzDM2xKFv42jK9lFes0UHbZTHzHs+HLePxMnYaaSND0Xt1
uAJlSmdLiScdTVe8Euu2L3o5N2TVgbnHSMmnqBVDVReUzIVXmBbeSJRXUCnbnyZ9cHCvaBnWZPQF
qoWu62xpiKLAMbcWlM6+EFPauLLXPfjvAZWO7T13fShzktekISJ5gqWcAcYNy74KwmcDuB4AkdJL
gYR93Thkbjk90QDYdp2YfBEH4/MC4xy6jqp5xZZzC3EYOtdLIPZFjfRr3XUBFwCZolKvdKZxi/Fi
hhNhDDoDxB5ZO5FNh9bMCsR/g9hRm6INWLRuPtRBhSS25pldWV+95s+F6JS1vfEGecPmQQjh0BDA
xIFU/qW2n5rpnvcLW5zWTGCxZnYtvgpaJTHeaETmPMJtnU/z7DByjHjM07NV+z+vjquOyLKBnqbB
J0q5c8nk1Om9d1TH1NjalREVKvzbhqCDSd03l2L/hw8zLd/KUHXed4xGn7mmtQdmal3XTmNIbJPa
1sUOUzZJBrPihz3D3/NET1Vy7bZOK6yny/ekwi5D0wXBfOhbLVCu3lG/UuH8daQjLHCFmI4fKzs0
6mBdwx9Ciy5GkOIOyXOoE7i5uMJ8qz2Tmau1EEI2DBU5pzb6BzQqj6yMZnclPhfS8QCJtBnOOeJ2
jrKCuKHzgv6mhAzSX6T8cGQr+GT0UkNME1W3qGQdyvhmmnL+Z9LE1gYxuYD6koPgRhXe/7eORWJQ
4l4vIUSkT4ciu4Ma1KELHaRDzot3rXePrZ+jz2Jhyaq3pAQ03Zz0ByOWaNSf9oHdJSQFSsu3K5t4
Ipan2iHRrdAwtCybGv0Mcy2nFWsRayUGuREv6KPKjn6dbs9YLguSvnGiiG5KPdvyJgNnAPSNL7ji
48qC3a068IN5Zdp9lrK4XmxC+e0zJDV4KgrBnRGK4JWxnetXtY9NDd2V/+Eapo7LS7t1B/Oou/8i
Y5FxvZLJBI1biazHvW+sxNBsaOHExSx/h6yGfpa7La/mE+lKFRb4gDq7tYh+rtf08+EV7BYYfcv+
cH8vi8O4/fl/RbhEDVdJClJHKwJd5aqtYdgoIhy+o0ZGC7tCB/TrPX7Pov8Bx5GonQLWqk8C2N+s
8QJuyA37UoqveSFSuaEtV6BnVjl59AkL4bZ+J5RrDRadlE90i/IHC+cbsHtl0/OOXB/OGtr5uUz9
JkVZjQdM5YWKTH2oiSrA3MkUqSmKxIo/oRixpghqvUFB6AUPsD0OeDEuUBroW97k8H2O8Z/Y/ed4
hyXA+O3ACnnK+xcqkU2N8C53nRa8HQ+09Ie3IqMUWnEbdWJ7QUqP+ZMK7muMlZ49qYMQ9+f7Lo1u
mmTObjVwprG1Mgjy7gt30MbPfUrbgFsHOjm5ZjsjDGNXpgKWgrdoSlmSUJQpvZ0AmBe15uGEQXn3
9xrYFgIwVTpVuWylYd6zELOJ6nrB88HTv66H4d6PVoZpzG0GEX3XG1LQJdfbZ3mBLENd6gTAA5yJ
ONYz8L1+/3yIN3K6SskNvQNk5ZMZIBujdBqCVOBCLFcWMAXsuLMQEab/0BwvsmkY3kp4Xwt7t7NC
jdY/gopJUvSC/zbmG7s5oSTQMh4OrhjPhH7nc/d4Zrr8Zo8vEsSusd3kJnrYPPJxSgBwYCll/XSn
8PPNS7o3fg4dMh0ZiMfuu6FLISsGT81vx+WTeJP6KebizZOpBrvBIL0ErxRkfR1H6j3mN6E/IzFM
waTbPwDWBFxLiZtYtEV+9ZD7ZJMEDDhVDzmqKJyHvKcFsN2FYcPn1d63kalL6HuyXBnBtHhiSQJC
CGhzK4/TDbDJWTQNMHcHHX7T5S1zW3+cpKF5a5cVwnxFJxCDC1JnASEvgF07o670kaUnsofuf8AO
sxeh94c5wa4aWdwOKXe5hklTc8M7H/HaSou+i90ZBT65PPZZGVuUUn18fCMDd1EEq4rWZqpKfTvc
ucCSr13rBQJu2J59m3e5lsuiDji53jFk7vSB2f4hI4EUJ1R0+LT/KMPHUgGe02g8UR7+lAoVk8Hp
4mLSTHY14LLN87TUtkHrcReUA8uKE/NSS4LQenzdjBT85sHK1uE6zPJT3ZHgP7/hYeBCTziQOwqn
Ld/zYYlmrQiVDMFSU2lTfsGgV/5dzc3RRGa5FIR0AyTlE1+IyWxBwwR3HedgX94cVdqqM6YQr3pM
ZYh2l2vNpfsHjD/Wvhri1JKbfqmfDvKquOir9t4W8jcgecGkwe7Xr0UQ8lLw95VosAFh7jxY+1Yj
Bbn6I3X5iv5beaWyLfcOI2l+tVpDeoG1XxNVcZLuj93I78BAefISswIS4rhOcv8T4DPrgirqurcj
IEX0Vyvw4atyJ4i96TynAWjBWJ9BPsG8eJvMD7wiqYkyM3xMVu3Wn1qzfy0yfO3OWAOazUUuypmS
eGYbhE6W+SXtdkLYLTN9sSigf+cVBf2CKet74PNNIDqcL5olTnnPM/VyKvPx1Vu04Ki+TtKhKRXa
OnYDWb7Y4C2CuPTKF/VweZaqLIaiyGh2WEtB89RQhBOnPYK5lV51JWKXvPt4k/uH3EyHJMNa5+iv
9+7adYhZ0ORL5gQEt6NsLi3k8jPb4EzkzAbJ95q+t0NIjOrEBU9ytiOf19HSZSJ1+RRe5gwkL5+d
OT+S1DI6LFDWQSpsA7FJ9doAihJ6vWFr7JG1OCGkqrJgNhaV3e7wo+YpunqcbZToKfgO3D2WFQK3
zqSqizgA53KQxYdMS5PrZtYSnASNwmElt3AslYwK98DWhamKB+uTb631EM+zkk/EZqxUcgrCGwey
OdgeBl3CQkMhsg/tGIvBhi3v93YuajsgvkGVbEGaEVWj6ERQHETYe6tNUXNRTryiCb5E4fw9l/IF
KqwQxTSwJWQeUM2q1OQRGv3L6yRPQrm7VWh7I8dlsN3zHM+VQ9YmbZoaDe1VRMHPD/SLBv0wdPjE
iTWWntwYndz4MqPKmzFhP9v+JEHAbH9vq8js9zXy/JzGrjGKgBb6kNXyaKIuDfxk9GwwmHv1C3Dm
75y6zR6+ZnDE1DIgPOSVqOQKZS7SflJYXJ/wwuDb0WznG6TTa4+/25iKhxHxHLj8xEfx+EQp7WDk
6nrxVQpREtXYLEwXzCB3iwf7nFHhsW8fHpwcoLAU/VctjWp6vJkLZRHeNVqA2WXQShEkx7AVNx4C
HR3lThJQ1YZStwDmBDmnQkwTyGTgPhAVsOULTSkJoWXRWJDwaHbYuM3000FjYwHwr8VOxXarc+jj
cSk3cX3QFB3agXZK8EFN51LJi66bI/e7F513+D0Dwcpgj9JvmEL5G4gUkoL3P6PtA8Efykk8P4jQ
IO/4SKVac/X5cJenp6bSd5wteOuLy8QjE74sK2v8/o7GklJCfe1dnE/7OKy/Jx4njIXkpP6d2Dt6
NYN/m/fmhPiVPosu40p0/tC+vVf+O4Jb8ZsteJDFFzq7SWjw+z7sj/gPWqiG2GW5UrP9wA4VwRAl
g+OEyVjagP1PIKkZs7extyAsBiFTpqJs0+X11tEgMqh0wtR6ta2CPzoXTvqii6Q23+UixX63cD7L
YUhWeAqBpoEXFjJfZinSWY+rUgOR3WhECsB2o+zBWXxYagApWgdro08kTIv/GnVSLx3phgUO91Gp
O6Mvyog4S5G27d39kxhNTgHaf5CzhmkrUy751E2wdDI296xbz+HAimzUokBmIUnSxqdGCLb/60Tk
hEI+LpUEYSgCOtFLlhMHHoSiQKiTJH5Rp3SEQrs0v89MmBaf7jj13aXMZ8VUqiY7g1jgt+ryspqD
h6laEEmutNOWQijhnhfK30Qi3hgrCR87lbXPMqoKkpXdYA4XNHbnDcXa31HRzhz8KI+DojR1cuiL
VbE9t0oemQo+MZInikgfEPZXe9Na/roYA16PlGcti2QY9EnOEB0mUa/HMptZ0cAsoYEpiIcXmCcE
5fGyZvOaFGhdr6fwmXlQUI/d5VReb2S8qLjuSVpo/rwwxQITp1mrmjRzjAmKHdnumdhHe2VRHoo5
7zQFz2aNeRccamYCW0COqtBC8WBoLTc42TH5IF2A8zZ4R4Dyc2RBDINAvVo/JONt1wSV+nP3ABd8
FtJL2pnmeZZqViVFlc9Tb2T9UCU48Bo60KTnHOK+rkP5Ba4LwpRlQRrsGA+dD0WLjKMLcAKZAM17
xRhWVN0uOV8x0DWS4rW+29BfLsKvzJsaamlAiDbPxMVF/qjACtvN9111IhjuGQ46kcCbCXruyns4
C+qdTc0g+zUdbVDaHZBPt0k6iF6nsAIRNuwThFEiLkD5vE9HnRPogLj2PT8MDi7UMt/HIu524XYW
6yNcfKzOClifa9re7W0MSgK340lTKeoxqhRMlyWOxtn+Q63CVBkeePQ0LQvYFRfIlsDmAFrYTe6B
Njvo4ZpiMdrLmX8OtailqJzJ3kD0+XlDJtGvTli1hgPlpAsjOru+8uBoGCGVz7XMVf6DsgF0vTz9
RWas+99kKgXv97rIQHh323ccwjlMoNfMp53s2LljAoj3qk5IC/b20fxiqYaj0ZwJGAak/cIKxOkl
qderhhIYbqzeGEcuiqkkYL1VA4wFHnGpheAeYHkAcTd7MfbLr1+OobXvjWwtRfNY6DUmYdQJB7BG
ELFgcYMN0OMKnH/pwwbxWhgDLOb1qkDlyvXaYdTyUwlaE/dyXc/bNR1J6yRRkBhYRaBrcKZoXtwY
x8XcshWfRhDrgV3dSFuBWUKSwCHym+sKN5d/KCwopHi7kUCRTMwyOaR9CM2TSpHvyG1HgAzpaxQO
g1dZ4axDwQ4YdWALuNs0R7WHrKuAa0zGT2X1/vwUrX84W0pqnKCrzZA8iGSHz+JUWyvH+7HW4gnC
vE05bsfhYDpEtdRDaTVF8T1QwPz/jl+wQChSEKX8RBAlUHID1SR48qyMSCnUAYVr/DcPq34v/0tO
JWxKbITzQebJkymZbEW5jXhUjRH+UahcQdQIjUS8sEmSImX5UEI0Gnd+cRG42RLjvYpwR3EFrlbb
551qEkiP6LGD8qTbcYx/TXRU6ENLnDVAtlrY9eL/Co1YOImeYZKfHWNeq492hkofHe4AUwEO7B6d
SwRVugtRqLk/X7akKMeRoVk0p2ZGs7ui3hMmJYcXTDC+o5f7MmoYhek+oKPiI/2+9ZK+IstbjiWw
3qjpJnjqwdJLuqWLn3t2TMjb4a/2SQqF/nMZTuXCn5BN+sVSWfqn868RissZHoO14RmSTcbtdUYs
5BIjrOhM57CJEsKsB4fVVaEBML2IQrpiEzcppMaAS0uwAmQjrGeAL/Bi2hr2GOeO7Vdpu+ZDSMQ0
TKpQyGyfpi3zyUDZG67UG8vXlDLIoEaC2CJbg8GtGDIpUuHWWmUrvukNs4los63OgzDcrzNyOzL8
jLJFXnZmTDRM/jA2tpMTgWU3z5nktM+PrpwCx+sMitFQ+bXFfJA92J5lLfslhExwyGg4rLUNMWo6
WP5jsZvwcuNx60eusCMy4yBt4zSgI4Z4o+Rc722XTwcoVh5H2pMFzSjYSEr+o8lauZ7fWn6eohdT
DKtLL84YEDcjc5K07Z87WexXfBDcNE6O8JJH98EeBz0PXKn/WSkmRrfpwOFaF5dwqku50XtFiaSB
Z7uNaWTjyfhZGCVAPRXFGy/APwcLH+6ovnHvViJqGVsb/oOxFAS1iJCdjjLKJD5Dk7c3a5JN8wS4
uNIdGYs/xB5qMHtmfpSPHQAUFhTWEMLSbONZMyW9e4wn9n4t1yw0Og+GTo2XKBu3QBiP6aCKR+7u
pv7REOZ1jYrfK6O48ZPioLNi9Kc7Wg9+Vg3VnS2JsRmk7W6zDGYFmE0daDyZKC5VL6QUNK0UHmga
0DlTTR4kRWaJq5ulE8RELUAqbFX7IOA+modh727p9TyW2p1OZzS+vD/PNXEw6WS47tpMtEeACeLD
D4do0a1n72zt+kMoPNWrNGubuTEpl+67m7KWnwxfLMzM/vyyhWkNxnydt7ZB8Rvf1wTcDNIoFMbR
ZBBzG3tFTbxnaAcIkYS3LAb8SjZlbzVCrlO4X0xeZUyo+CiDph9uMTo4sXQLE6/hf9Mv3/Dw/3qo
15V+ZDeqcjSwnk+kzBNHUHqo012HYxFtmZTnrCpOqneXwd4Mk/c1BRjSNfmBvIEh/GFEX/VlOlrm
QmDGsiD1yHoDRd2Sf9B69AqgNO7jQzStok7GVXm1hre6QK6F7NFcNmv+zxTqlqLmOktrX0Q09fdF
ekZmEGPcS8giAEDnSRQAdtXZ0pLf5fqUVtoV95vrgkXwhxv2RyuQdxu++Xg8MgCXQtCa76XNTdXA
f7nK2N7O7zJNjahuuUSu6C2ShF9kJVfQYfOYki+YOQqlINzoM3ZbL6M1R5vUpSYuDGNM7jn9/WMg
s2sTRjKERULj4N4Z9K1H0k5NurEcks44BphVNSsDEsNoy/ll0cUwuMoVo6SXi+G6pJx3L9YPuh9S
TyedtyYjTNNF55o4O4I8ZJFuH7T03cONAZDYC/AedqYbk3KlbMLyHukTJBa0ctVRazy2dM6Ve5mr
A10ozcUurwiD71yEe1xctNP96sdidLYRKOK0yfLcwA0Z0qRnzPwEc1NEj3UC17ShzaDLKi/fvIU8
ZY/ZryoIM/9ADrt5y3QywJo0zXGzIqDMe6Xs5oNP1/7d5ubl6g3AKTFKSDDrdywkLd2hgDwxdlmr
ZqjJZppMbc7+vHVm9rkJwu86p2Iu21fp2VWO964E3j5m82whzSEMTO0Rk4IR/gQE8e0JTa/GmyIx
OqD/JFyFkihLXH8eaApGzFzy150j3N2fXDFkNSHxIcxjcAOje/kCQoS6Qc/N7ah7jECiffB1CEOr
bf/bmN07VXnSowFSuVqW47sbMCzH3pPe6nG8tIGosTyYjKyVxaRldsbYQNkRQnhy+W9hzosAuzRU
6dzVgUyHqIig7SsRTX0exrySICMhiL40B+NAmiYshUlLFFnVQ/yittQhHQbfGVUF+SbskIBjdu3H
D4/nkvd0HjGf8sm1a2+Ez+jdzV8fM2iOOSYM/u6MSGXXNNGzzloaki6pUW5XTn5PsZCoqGFQC3nP
AjKupZqQ18sqga64et7s70xg2xsDAY18SYdVEOMVrJgOEnLE23nk7nwQPvg1DZZSRxUcdQbjTymo
iLK00ia/0Ls3GHD91iOI0lo7sV4PvW7UW3acm8zKv0/CXqTYpKaxFclI6sFzbCAq3TKnRUoPddFW
8/8+xw18NShTSkHHl2NIOnHa/H2sYWu9rbqO4p/fI45N0aTopXyf1CdIwjin3Z2VXZutT7ovuNti
Ex91Rlb20+tpR5LYq1lclCb6+BXg4J0P7Fauu4b1bY0cqRmY5U883CaEUzzsMywzBdR4vjH1Sd4q
VFJMAR3dOiTM+ZB/CIqfDZzAG/8lk61LYTLUL/FWx4wmb2ZBD0eJeOEz1u8wu5FSY11HURAzSagc
DeAtQiXdVSiBuy/r/yLFGFNX1CDbbuUJan593c1aIP7Ui64nD2dCSib0f0uxXyh88c0JmXVvi/pJ
G34hggkkGYH5KkwXLy7VAOkeM9mSA2UlXNbEtR60z4tD3A0Euh4hHhiR78ym1Jf9u3XdoRxoDFqp
jr4HzGngY1lLhRjhvA0CV1R+aoV2GMJXbKYrf0NpozHqCht1SVmajXBT/p/pOArEH6AGwaJusW0h
LytCsbaFlf63M6jozpMh8Me0sKhbd+etmjQXnbec4MDwc8eTH5Donw975JjgXEYHFZICbycJ0jBq
Nc70tessKc6Syc7CJGt6CLH5WkpJTzEjpayft8NAOeLtDRkC4tP5mcsmMJo6uWzKi1BsqLpR6Pyp
40CcgiSoReIFcIed/9lfujrEJk9E7iCB1E44m5HXn7A5S7svivSj0xgOq1LqmpFnTCToHv6HKs9m
gbYNTCzCTziwGcU96wgwEh9lx2PcOlbbuyP72Go+fnBeXOPPNQc4BDHXJCz/SYEJl3EMVbyvkUHu
zBratnSTsDAGxhrtdVN8rO7V49BzH3TEjPq7vXIeQGISWtfPLm0HArCnFswsVi9vP87qRAtOLS36
ivffw3FDHd1CerLA4Yzp1H5qz1oYcuNePpRHZMr4SDUB02tECnUJAMVgz9OU4iHaiAp5q2Bxgf3z
WsoEwILKeaf6Cxdj8UVJws0sRbwDQe0JeVsDEW2MBq7sj2vOzxGLuQ8cZvyAJ/usVbGcHoQcaFRC
aGvo5P8lgLs1NLrru5Mp4jNce4IqeXpHFh4arWsNafkf2uqApS7InceIpVKXS0Bt/mt/74fTebLg
XE8G4EyIIdJ2CE/XaI4XOa9bY4ox2s+ZPh77Q+P54BzeJKQbtvzkfUMw+pMSkKJpqhjZDxTt/UMa
ffNO2G+73bUzhT5nXROoNMIzLNKJUUsR0f/SA855d8QjYQ/kWiHsPKmrgTBv2lLA3+NgINeVuvlF
BFIk3GAmQBRYQFgIjQtK0Vhq1FHeVAdqaxSIv/+hLNa/XqjvGUQCwIqVjyxyu2bZRu7Nzs/v0qRD
U3iAZ/kcTHg5LrITyUHb0/jCpk/3UWLVnq7gCCmVq02DE0mP+ERgqcdtCJUHhZhHRn5T7fuIb/ok
K8EotszIX8IQM2LW0qJRCUBMr2TLQoWmqx+dZfzsBs30+eHQloERZXCsQGMBMIrQWwNaK2ZHakwh
5MpthXtxP7nQulYmrE+ULMJe3VDLq774Dx5ZLAvOWXsLl2KV/OSyOLWJIcYyZCBBZlgINLb5Y0A4
9gWsVskm2av6+YSL92XCQx0Ve0XuTZI6SHIk2o3uueyInVV1f830RJXYoLZms0/QYWVPmJkpxWkC
D8krEEi1ziPCHFTZtFn/ZmiuBVpjX/uj2n/HEdVZsII0nCabxxO9s1YpyME1XQOQIfMieDPYcH3J
UJaZJGBE2/r+am5WUmr43WfCPCoptmQ/uEmEzpbed1AVAxJMTUpNyNbeJ2iRHBPGgqt/+zM1Y8WL
5qEgO34SykBcWaioTZxz6uzBbQ1WcICQIBZR0cvGl8nh7tHvUMMs1XjSg5kxiyzV5GfoHWZ9Oveu
P+VXvGbJE21KWWTBhDHHugj91s3SrzFUAGRzGxKjNgpXdxrtbIJtpPK8+Bv2BoHg9JbLAzt6BDR9
Pr2myMS1zvwS6F8/hJE/uIuVV6KCLbmj7Z5dMZO3jGputfNG55aQ5VDvpA3Nfjel6b5xZjnoZdKU
sWOeTxkGwXyMAYA29661bV4ygiRDrlhDTyY3vRqRGcWAOHtFqJhlU0xDwXktukrHPCq9WvmJWuoM
j4DlnN2mi0cOyXGmyeQ/532tSebcS3KPc8wWV1d5/7rsd9DVyd0m10iS3AnSeGEnW97buSP4LJ9C
Hj0mkK0R9NMvto5Omlv2RQz2WcSgR6eMunlW05pmfCmDlIwktd6AA9vR7z/45ZlM+nEo6GDdhsLl
vCng0t1n9nQ1fb54YI7Qg3xaHFf5YZLk0axUF8z+hucRqw0WmMP4o5y0kOSdQc4hyRlB4ND6VSD7
ahFWRmmJlKKeUpK6AUhhOacXzRcieQITqVcGPwsz1A3dbQV+M9kzoWAPbOEZyhFRONXL4gL7klzG
WuHZKOZqlVZ2xq9TmdqnTzltvvk2TLnj3UvP4aPNd1zprI4X8SfYrBklC89RCtzZYoopedXb9hnn
jqciHGI8I5l1WEh0s82r+lLjkiiCr7A7Bo3NguzFjyOtqxzCVSM8I5dbqef/Olj0L6EDPKaBVagn
LLxkYZaupQw1PquM0uj2wpO8/N1tBUFHpBGhzE/t7UiNCnvK58emtMgUnQGSMc8gcHTPMhONFxSX
jb8QEqCgJKEDizcpc5DqQ/0v8hW+6eePCu2bvQunTLn6hm81sKzv2UrGYa/+y5RH35B180HWhDS1
uNWa2HQqfCPIQzKgr7c7Td6rBxz/s9kPawiwVxYongHy2uF4mwb8u/lRTmNKHppVXkTYk3ra8oae
no6Vnj1JXUxSUe+yf9fTPJmy5ufIrOSQ4uCd/Lr1wSUNxeSw4MRNmAd7dGJ+EnXS1h+5Qh9PrtF2
DP0dBpINL5TC4XHkgQ+SPw46caPuVTcpSINPfhD/KMEKo5v3okVOIf9ulNGhALmPAib9nSMWEOeW
9fwXayPy5vLvQ/LT82FGOO2zHxdqfpGSA06QvR4wGvGz6lb4jt2/kutmK7fSfrbRZ1VJmqOILhz7
WghKalB5zOE+pNhwZP5AFzgFK9+WcpO3I/mFEyIHUTOampjxi5EHh+iFJohs/63Ezt/2fdVy3mQf
3JIkL18UQdC0Pv/g+yWkahl4ImfMZ2+zDGHhuyFKz6YCB4DyP8S73cfh0GawOHRrvU0mDfe1FBp8
bm8jwvMfAA0NGPwmG/2bGWkLj12+zPp34XZ1z5IJgjCvH7sqg6U48lVNt4vDUbLKV/xJMBpu9qXP
SLpkuwPg0pznJX4nRgtWmvPdis5nCsltI6MJU/xxEXgCCn+AGAeZ6TuWezPpn3QO8yGtMFl55ydU
D5jFjtUwC4f0zQYxjCPI3VVVujlp3nuUMPIdJPpCwEoJIGoErr6altLoouC5yVrb+MjxHuMDtEIH
6e5w8W6+EblKx2y3Keq/dBFds/5deTUQuKqtzE/iPNxrA6F3CkTmMIhIQWncb5PeXo7WTy+0BJJ9
KyDoXr/1Fra3HWC36rKF3TsxN+nS3yI2/8Aa8AM4//CgCm/Jq/NY8bpW7B9nY1pkN09D0iTvOrrs
QPrCivNS5TVLLEd9Pz1hsGUwC/1vlsJlmZL+GxGUQq6Y3IGAY5wMeTxgIOVDF320cfoiwU1c1qYh
fcJyyN/zDpJCSCBIcs/ARckYDqzd7SiMpz2ZZh0Uyht2C+0zUvFHYnPxD+ZYoT5aH/gp3fO1UrH+
pQBKewHMc1IABWtBTJVb0X7lKN/PR5L8jOLXf8XYUURAK9lDGbhlAnpV7Rtxr8voyge/KBimeiNg
LDsiqnslBZicw5UmtI8+sE0UgwR+cHwrnCL4sSEzCBEOGEc/+YsOSwi4weugW3evHaiLTz49SF+5
zJYBR55FUOyy20eyioGYlDzcsmiX2OBU9HeII2hf31RFh5kvsoaBt3B77mXrVE1C7vM61LvfyNaf
R94kCzEQ5FduHx2nnWBdW0lNsdmNIUCWRIehGpgsgJBjNqrv4uVsLCoRK2ct/Fq3aHlxrIJIP4Jb
yFTSPbhhG8ttpPdBu0qtu/k0xCb4bhVy1YLzuESSsd/FYQncpyLr3zIAEn9cX0bnoZj0Ess8kje2
0JeXxSgN0IMfz2BS4dMHzkLq2tl2z32+dP6YKQ/8JA7HNEuKLjeRm7Z4n8tAh9zOqGG8iRt+cu8Y
VvVCSFLmQQtDdMeq5kBIMDiAZyv9nGPm2CZoZSLquBPsH3FLZ++NYTnOndWZp5prGp8S6DbsHpTX
0g0cONBW8BPFRK/a6uJM2PeXRIQVheoYsL8PYDA5KM7MKXF2eOPmP2MtpK1yyyAXKDrzCIBH9FxW
WJMkezqZKFGNqar7uy2cTDMr9mW7XWXxrzDRUxP830upRWH45rPQOG/goN55oUAoucNgGG1jtY3t
nfaRLcY8QY3OfL6BNBs21Oov4/Ccw+mvOzQjJG4Ohk/0YnlFOXeSkR1g5G9wnPBc7LYVj5nXoc3s
AXoMv7k/s73OCGIuUR4uQ0e4GbN8xCgJ6PwMACysnqFVx0X45rh7Rc6NC/pZbv0YtEqt/nXEt+Bs
Fmnbx9pdTpOCewPp/OIxSv3dqL1sTG2d6FYwZaLR88cxDXe8Ratvwh249gdN1C8jWghesOqf0PgJ
Xxt6Nj8UbD70tBowRhVf2dBu4aHWuzE8HTiDDDH7uDyeJUwyIf+tGON6TreOBh8ajEcpKHSMwtzL
PUd3tSTBJIcGCVSbUB3yO93gjZ9OhaerbiZKXpiTSFvxhlVufS5rrSCfmD7zls13GNkZoZii3D1q
8B65JND/A0SHDr5QrSiUJ0RyOjxd7Z1bPQOlk6XWIY8FGgY0OWP6kNt8JTIKUNCV8IoZuXzPSAIl
JXj1/T5+laA/chXra0kNIbZTAfaHaEpYddVBvr2bUvCFUTjUG7l5yyidIcnaGop/v5S61E8oBjEA
9fNM9QAV1ySZugAtnyO8lp66X2m83d51qqyO3X00rBzlCvZIgDZvU5IQicf91oboH3DaFYggS6m5
OgG7IP+d9sQIVFuRsRrc/zWaasfSXNlHkECHGFyM6PRvtABz3LtswJ8o0pnFaQ6W+HqiTmnFrfT/
KtjW4B0nN8+UKG+clcWn4SpB/Do7fJuB405tR3/yoKaFWYgfE3gRXXvjBivmn0tIydZXLhpIlEEb
lbtyAMqRnmPDXnpGe25RmZCg5X+zpEj6b712mnODJkni81ysxORwhrODRkEEt80S8POg+WBgvuog
vxZkyDgZLkFdvCq5xHKXBCTxKk+D8S+D8WGVX0qaMDXxEYft2cxlP/Goe81YUV0blwXfC3Od+kUr
3zWf0IG2GjOFcQX8CEPT9y25pFt0OFMjVf8GwjyMlnP7wnkyEyErdfNjM0Ww8t05YN5D8s5a+IOn
eiO7z+wWPenasHtyNRIjAVvcCo+OQPuXzPQ5psupsI3umMFyMCLZ04SvcdOhTVex01bcySRnNlor
PzI9apMxJ32cOKrJJd75g+04Mg1YgFgh0dsCDEpAJdk+33692V3zg5JjF9czB44hMs+KW1wWjyn+
gKls+hZAtavvRRzOzPjApOPI1K1QrWN1XsYfNsnYn+U+frJOayC1ClJusSe/8jUq1nYGxfzqoBqn
jhnMt0Je57Jn5PBLX0kF+HmrIGZTNE9CNK+R+R5hYMcg+5CTRibvRe9QgcQv8CCkeqpWEdK9s+n+
e00Bskg0rNnYJVJoWh/vNuCAUc2b4rYfz9tizSH1UUT0VCyfGItWheorv2m2eYS8yh5Xde+q4PvW
0Fxiibzw/Q/5bS7aIGEbIAxD2KT71G4J3/lO6cyHA00q7zH7sj5tDOYrllIbVyJQJ+DJCZppUzne
hzc1F/TQf+hudk78VLCFDV0v3uYa96e1KFYH2X6Zpge6qxdvERy2HIn5ImW5KsrZMHiF9AE8pz3T
ia/RKht5hbRk05elsMSJbRuR4HzEnGM9L2Jj1Y0AiGmFXoLBPb5hBgQzqzT+xy2wRSu83bKnQksf
Gl3icn0JStl4cW4SMfChWAWRDL5RrZo+kZlPwtbX21u+fkAkF399KLzsedMfsm05px4OSTFtb/Ej
tF+TkD3Xb2lwQkeFZ0hadsxo7IGrO5HeOaYM28i6rYpZttiWVxUfVaUdfiyuDyNGu/6nLy9mq4rx
tiLcsXxHGAhHqS03g94LQccgnrgStjqEBz4pBZo4fhoRNMYsSY8Dm86liep0hOkBnqZr3InF5YRD
sjoyHn18li4aslvRNgcJaXDMfjhoQTO7sjFrMA/b4KyPMU1Fq4N7GrQOo8wgPechJ/wFziNTIgQ7
TmwTO51eZ2+D6hZwNXvNjrtDO95qsSk2wMGpchBoh4BiXcfbaJgdoohUZuMHRh9wwj3K8xnzdCRC
oZBSOu3dJd4lZTaNkdIQzR2XVDkiojlVt+xlth7i2PmEsLeeLwbOsZIO8srPoRY7OKbcc6nqFXXy
JNuZvecrmyIDczAOvpFdhd6+obgzD9SOAyGeyIk+ZxFbyyoruZgmPqxDlMIpZlh1C8USeNx9cbBS
g721DTNLtBRaFDgzUBISmMikl4IvJrt9ikYAKg8CHq52Uz61y1hmUzam9lZb78ANurmI8Q5fcddo
1Kef/klLxgKTd0+OQwbvx9XH5LUgIsq/9b3Jml8gOjIPfAQF/jBB5TomAC33uXEDZ/8q1g8Q+y83
AIHp2x5LIs0K1fPMt0LD4M7YdzsWA30nfHYBo3wr1J+ij1xMSLDM/aS7yENtysn7chlkR3joSutn
F4+fY2FkayHQN8RKBfA0tGoPqr3ouj7r1kKy3KEtePJmEiw7D48vvyjyOVi45IhUEsIbgXNlGhTu
WN8+J92DWLfI5Xfsp0AiK6EpdBHb0Vryy4ETQarX2vuKYpOly2psqwC6nFGuBKbeGKnuexWz2+u0
099eF+MKVk+MIhOEwUVZTuM1MTt/9RTX2zUQOKZ89eMinRS9C2b7m3u4fOpI9u4nG8cq275byfgL
94ujEvIFP/LL0gGOldDzmkSMK4A446Y6JW6Z6ptrdPUcjMlmckC9iPJj/D141MIFbuHBofRDmqbL
FhmtDudHV8Wq9Wt1TsufYDif+HqdIXytoOq0r1pdQMGODwm7wS1qjGmxEHI5/8vQQzADZCbYGwwD
mLtteDHshb9du9klLUdY/BP/ecSjb3XhREer4d2Ow8ARepxyyVeDHHSGeCUjSXo5AdWsB+T2caV9
XZThDP+3bMTXoE3hFM0aMmKFb+0AZfKktJsbTBJKBGCCRA/dDVfXGyeoBTv1QPmOYRrc2GgAzSUn
2xeYc3AcXfeaz5a/2jiBX+PlMG+8DF52oL65/zTtEmlFk8LxtEeL50OO+on2kcwnnDpWMHt3zFfF
QH5fU5B0zbx+Sykrik+9tgTYZnmDbzPZ+IlsN6VmUkGywNGXVr2jicUlTT1XMB4cE1RlmCNes6qv
Thb7J9m3GG3BsE7DGSnRlQgckE3AKDBfjxE9ShqI9PDudU7mq7NatXFzwLV8Wadz7CD9cXnHRW87
yWAHh9140IKDqVwQhm2gJc6q7V2i0QBdLe3IHDUyMk/s53t3+jgUHxqmWxMn39kqHQa1nu7dNxKK
iUzcgELD+9HxILCnJvaLILdBWAy/5gPO772H0NMrpg56Q2Sr3F2Vc8WfvX1DIm29Ju2jAl18xgqK
ZCQUCnocILM4QuzGd2zgXOnoeFEMn3L1WEYe4XsPbSQxGgqrCryttQ+3qmefqbegz+Iw3j/1kthz
aSjc0PEsZ7qrboz/zZ0+dKDlT2plusJgKR4nAH4LgMXWyBd7+K6XFNSGbXmMes/ES1CiP7qTPeoU
g2hNoq8jMKcb3Nqy5gqZfPsS+Um6i/ROVOvXr9PymtRR2S6a3RKB2EAvlK0r3O6vfgHaR5ZWCijC
kJBSFCAgvsXFb/5sHThwo5HljrdS45wcx0JWtJJ8H421IcujmK4w79eLEAMu3X1XT14Q3PFAU8hs
nNmDEWLAZ6Wgk/ZDMjUQSiXpWJMn6z2vMP2Z47w56B64PjE3jdsZQ1Eyhj2xUHpj7XW6cq6rgSQ3
uVJr/+R8yK0ipoQX57mfe8LO4PdAe2Q3Su+buSZR8mu+NwF/39zqH9QYqQUtaVFyfRscVK+p4MXU
zFFR8MOEMeYguhrFqIS2YDRhVvtnxHQqXtMjtjvzHkAoAL1Hm+YngOjoyB9rPWhcsUTp9bUTMR8u
4/eZC5xL2ZYY+P4U5yY3extlfWoccyaA6bmW1+bE+RInWv4tNRjs7YtFGOJ39ln9IAohvhJgvCod
SwvhJoxQh1jKCWgis4qQk2QEB7EDzAXkno4RA47h0yK5/e47OcjDbPizRpVrl3LWzEp0IGwEua41
Vv4O7XkXtM01QZa7QsNQ/97pTqeEdJEw2vuxA6+oxKMmBn/IORlyKyAsrH94haNF3iw9nqHYpfm5
zEDA9YhSOlefWv/SskUwEe6NJcM44S0eOSA4j7gBxv5eiRaNwO9ra4RyRXbMduIXO96yZbmLm9w2
fzWy+fr7DjC0qJLlxXd+a8fOsehHXdhXF/AUgoMaAJuKq4FSY+1IVY3ows5EE7W+BPRkRDTfp+an
kfVsuNp6TF/wS7Rq+FLwCzaKBEiXukxtqbHCtMPLgmJq3LjFO1qIJqI8YGrXhgbG49LpV0tODmed
ypFWzpMLt8y71F5abLF/je62yJfVgnUex3OxLyX4ZcBfSCBXy65ugN95qRnKTOsF6VIFBjqOaIkb
V9xeFKHM7K/Yt4HMbC5sp+qeaQzcDWzsTNgwYCn9CF8EfXTlJU7dWa6kUoF2ix+etEXNjesRfLnN
y7m6JJTSS2jjN6QSPR9TrZoRLdRBSRD+3C2A/IHslJsxN1ykdgR80pWWcc1Kevyf6PqGFvwaDxDN
o4xBbdtGYdSWJJeCKo2RpyVo6311Hfe+u7e44XoK4hmVSNx8FY0es6LA02lrsIZ6Hby5vn2Q0aqw
wHP1h74Ai/PJxrhxhC2cT7V1NmwzehjKpdwyNS0r4a5YP7DCVdAkempXbzrxehdEpc584c5cIRcx
CMHHdr8L5Jk2MRHqswDCVmunRwx4VpBb2ADpyY0HfS2kGf5j1q+op8RAoHk65ywIEsgdQG29cDJB
s9iXVHxqf0QC05cQCWAp4JO79nxjZQek2tdvqZkDPBiT2z6bM8sjfzwS3p6yXbwaiJ90xrq+jVII
aDqpfMEFe3VMGBxLOYRWcF5V4PJwQmQ4P6/UqIrsT+rsXIks7RwDjgZSNPAvYMXeryLt3BK5xUkW
wkaqViSVB1/2OOL/oMQpAFVaW8SgikHyAfbrwiBuTQtSWKEUJtZzvWZArAzOU771SEFAjb/pTATJ
dWQ1xxCaszS9OLgHrahK98kizROJdVAfwJUAX/RSRcQ1Xs1d2rYcXluUdGOlLLLmv37OMf/xGmLA
tjk17UGkcWzCeJkaXCZh71uFFom0LmF/JFnoQ4p2LykVzaG5UVF1HT4w3uDVCjXw6YbjYaPa0N/p
vXIivSA38Rx+IsXqZ+Wb+6XFulPevhbCcI5FYfqZpRhkVWuoQ7fev5pQAzf1lvKWxs9taibU9aHV
RpCxGd+P5lFUTUc8sCAk3Vmqqn0lTWyahL1eeU0X7S/QmjcJsEqArrtuQStqKoPJzFTNSx7b9vC0
Prfm3qS0eZBgevUZjx+uEAMDgJc05PXXb4Tpe7nVY0pNv5jixf4ex2dkdISiShjKT2rBNj+G628V
pYnXWIh4IPSgyjkaRH7ZIluSi2UBHyNjO4v58RduQLVoNnzmxFpswZq0oN7pLf7aBS9FHvVy5J22
p+PnKGJ8rh7i2++CSJKstW1uojIqsMsfh1xTpdS0q7gUQCXBEm0HVowSdBlbss3iCWkech9qK25j
BlRxIBiLEm1qXIlmDS5pjMQCadmJkFzctY0VJffAzgv2qgD9JnLWsu10JSbA5qa9EQGFQovZyrq1
eJIKJyorOOkLicTRha1zfRzkwa8ZJl7SiSx1DWxlQNWiqf0tW+ztdjkuXb9My48AgGOLlgVoCUOz
acD2ixs4cMjTkuKPO2hvfXQ44RXuS02s8+OdAaDnY/nNORkii8xmT2cvQpi3XIaXbhXWbcnQp9CS
8NOKSjSpL2thb/yNtWNFV9jJmP70AcFRwdlEXMKfdeCtMxmZJq9PwA7z1PUeTFwi6784KVrAapf5
5k3EYzidHNa4WqN8+CqJoT5rwm4gspdx2hY4xlflLYEXxmXdSkmMkz9d0D3iNygrPxF8SbatTEZs
Xb9gyIkzodyZ1kw1+KpERNWFP3a73OL3E47yep4Wrolk1t+IJaTeikKNL9DUEj41pRZMt2RUCsRs
jd6CJAiBWm+TkNYrtsWVYaW+N70Wy6rx2u/1E203AdWwr+48L2fc4slqbdIpXRH454tx2va2XLKS
C5BGKJvwTNlC1+lw+uUqt71GGHcMW5a0R4FwA92Mf3t/y3LBKiM/uyjsQzwdkA3mrGtUxjEURLch
4eC4ehH+GGPgDQcnTrKETjPsA51AyNr8N2O2MyprjJA0DlyHi9EBNtr/Ug7RU7TKWqbw/skSbmlp
998qKt/IiqAdQl0EnMrGYNziIux0sjEvPmdVBJ+v3oZkC+3hpsdKvo92NU5vkMwWR3rYP0iQoFaY
pSzrkjXyqrHMqeNC1YfO12JF11ko/sMo0Hhsgj/L2PcCtgp6NQPbi6NW45ozsYRT7xaQrXqrJLjj
qpSM+AsLrcaqKwUmLK5fSe79KV0ztg6PMBbAX+L3cokBmqgVVfb8cime0NV7IWq5JRb5Y4LiBFwv
bujKxBA4+iuPQRUVhlYPjBsHuiToWZeNmWRC7X9ycD9QptvQaEZfioYEGcMsA50u4CdVju/VxBv8
AOqCQCxB7Sjpj4qUpahrONL4F+CyC2KUyIADOyXCtbBekN3qyDX7YvwVA4H8/nG068dltupORsoj
YyGbg3ppciJ+y1hZcDKLiXaq/OiGHDK6bgXKAnv4jGOrJgTIrDo1FcgP60kmN4UpkjqsmCx7A+WJ
PTD6vq5Jg7LoaDzJXoPiuSpisD1SpRY02lowbZIhgprVh9wKI0AKwKYIYYMqEiPD6DhisK8C90xm
QgQndQa45QJ9OLUfkedikdEFCWIZo6+WshIx2DminSypowvgBloMOHnrLBr06tu9QM7PK+wOWkig
OzFRBVe9uVPE5rPJe4/Sz8bF+5EANUVY2Vh3ojZjchqvZDhBKm4XPOUHsawqmQK6FfZxs5k4E9ng
66NH/wqcm3OruGDcZCQ4gDL7j5hTxdtSR7olzEC1JxefJ460i3Xv++SCbNl3Rz/WXuDp5Q10RAxg
fx145IWjUa+hVcMFEPtg1fEpaymRSOAbbT0xWVq+DQjeUmqcuI9Z7rJgGrD5n3Lq6ATfSXO4SooT
OD13CTzQVehA1Y3+2MhD/QMHgl/K3l+kyNSMLw45ZjLqSNgGuvhh9mA1QJCRFMX/NURp2ZOCfmNr
r30AOG6GE/WY2VkrUfeKK3imLtoStKEjCHUKwFfJATgBQgFhgHZEk5caa4JTtW06YrVPUTyTUFNu
XWYvN10Fff2Rzjkuf6ISLUvezy8aBvT4FX236zztAGVgnk+OM0KVPW+cLFhnU2VY9JQz3dbq3nUH
w4X9CwnVYjgfa/B0msYIFGAwW5i47qnFMWYoeT8bpMkfG6zCey+pIxRwDq+/xUQI2i3r2FqBTea1
EenADrUKDrZPBjNoxlHzbQq7MK5Ny/qUkrxZJCh/yIikNtUozpVyjEHUIA1ABJL/tPz0SkmsCSYl
nC58lToF7t9v5cuNfjMXazFIYKQwfK354U+JfXwEHPqDDMeHcYLMxxjCuuoNwYTIbAKuXLkJ/K1Q
p/X+/l6IcsLFN9t5LUIYToAyxkewoFCX3m66GdPfI+PAMma0+OU8zD9zFbNNW5CLLf3gp+7XjBP/
qNiopsRtuFAAd+IyTcleOfwbaGDZvdvPknIxkbxPygbZJlVlY2hFnqdaum/gXQKPpIfnqYQ3CI9Q
7R0L3uUG0nzmDtYEoI8yGO0Y6KOz7D2Gk7/2RlsRjIKpN90yPIOPMHX00uFtZH1UcRvUDBpky+6Q
xyyjnHdJ/+g5PnNzHwXDfTtpRZHQGSmja/Dx1p/o2zK63Hmx2Dy8w1QkzSXO+6b+cy+NA57W/e8u
5pOe3tXilpWWH723MwuL7ieHrjQ95EyPTLxda71JioZwCAXphdyafbres+VFjcQDhP6J2pKbUea/
qEHeFNEIv8EKFhuBB5So3XOdrIOpLgc1UxPvEj4d9DE6gffahcuSffXh+3YB+g6ru5UXiUtZ3baT
uLcWETiFRnb/Yvg6pL/ud5yfV3TpSyj3ClVFly4YTql1uRzhxYqet0Ft50gVoT2qYY/NG+A4Tz07
abN30aEqL4oA8IdwySGv3133GnI0ggfXMt5tu2dBfF+KlHIrUCqt6kw5O5pmTpc3mPWBdL7aKq7h
fMx2Rt3GiikRTLPa9XgvoOVYA/a8UkwnzPL+pcB088RVWRZyoSQsmAhzjNhsB1CrzLwlPNJ6F2oR
2p3oHXWvLvbdmhsDMIgmj/VHfQTDfa8jHGDAKJMhy88WkkXdX3ZYeUa5L1QjVrRwTJdzuhY7AiT5
kzWVR2ngkh9jj4S7yw5bWNgtX5Nj9NRl7kJxZPfq3J83aP4CL0zsa4H4z4afpAzl0NCa9hwkwZFg
BuI7i1FUrTEztmd7fvlyIb+VZEfSot0invrxTXOEU84Wg00joYQXMtBKQl4ACigK+422g7v0y0mZ
la3jmw9WE62S5HiG5sgTrBrh5N3VQqjU4xFiFYAGZ6D7nJ4vmsQfmIHqH48NxuroPNYEy7mdybom
J4KkBcHQjAO9jW15lrZHil7hdivL2IvWlr6zQ6W8zcxOGZ/suuFZEeLtpfGVOB5Uo5RlFwrzoetE
ecWdbqAr7cjQJj5nEQyvA5JDGEj4KxCUHzZJ9UZiPCwX5vJbly3O6xWW5BRtTutOXR4mqYcSOu4/
fcbkpkauT3QrNNw45IO/E/wWrPU+UpUUkHLSRuymex2eShfZYlISqltozj5sC0GBQrVdilylUChh
crc2/Y4b7U1kQD1t4uLqZF4GVsETsP3pCOAYUWolnNfNY6L5eu3xR4Tw3BbmpXZhuS4yG0PiTBxE
9Ck8SDm0RIWQxyZmk+lzvPE77oKAjRT0GyCSmOsIxSWXT8W4bJfvoO6BVvnNnylX6QqjBNO8FSSj
wg+yJ9f/4VjUcg7z62uqYEcZC5hnF9PoyAUW2eg++Tv75ff1OPYUxMmrYGLZC/3Oryw78N4wqUAN
mUzqJtgYYq3L2ZnIGP5KyOmAhpGRS06TD2l5sZfMCxnkiiHhZRyQJBedCny749qbAqnOrbgRNfLE
TddcRuUTlbFxyDngkieHp2rY2gFx550iMKg1tTXx9roCI+PfAisthrhLYZkRpBC7pOrfOsUWcU22
6ktJ75ncARsF0BO4hdfpxcwNWuQNe2vmbEBeaAYjhaAfXB3Mr0ilyyzksBJHzHAa6lcX1CC/6yau
goq/L63VoRwxMdVsmjk/q1nc/rm+F15kDQJpM/qZZcVTpU6Nm2OQBjehz6j99G5NGaYEw1YHO7yN
dKRtf8EOS5sAdEAn8cwvIPcEXd7tzh3csfC396Q0MvNbSuSqznFk0Qo750lle83hlzk4QoaTRYoP
D8QOKrExgPaa6uizkpZT6K3UyZxyLeV8sLYpwGtdsbg2VJAHHhO5bVslx1JKyiRj569cSAn/YExw
uN4s6QixnVh8e1OyH+yln6GLkQBWRRey+cfFBlA4x9+/GYi18M933+58RSVhXPFiUEUuff2ZhX0L
hjAmXVofuB6306tKO02ho0W9jxg8gHqU4K5cUM1CUi/QgdCTiZQkR7xupTAN4/FLeOVfFv6GKtGS
oUSbQumMwf1mB1DWfjpoFTFbwNYoXGLm0k0DtPogIiNCtOheQvxTOBBgMF+S9fhsFxR9H77ONB9m
SMm/zmf0Pw6Ao2i6+x9hWDh8bdJJkTWTc8s7s9V07jOsDByvN/GRahEgqjXvWszDouCyuPFxMcR8
7mxkj/xlKD3huAOLGMEgLgsbBTX/zy6vam0Qa0LjXzby6mPppC4w3sclwATsqIdLFTY6WW4yY/vj
1ZeBe4aWFCiV3AmQzNxDU4VcQLNbxHOZbsrsEEo4BIJqomOl+scKAwftUAV/JjvMR1iRCCq4ImBr
yI4ntM1a+dLMdPZtrzxftaII3pnAzHVRxkks9Zzz5TLTIbQETylzNFMmwQBsff9jKgk6cYEFnK/n
puLmIigsH3IaEcXU9Qsev3mXidBglx6owj4IEIfwB3wf2zpFUN14Tt+PoqtVPBdFlyVWFM69G6I8
TSI9ZP1E1Bqrd/36PHj0dOKDHkPsrni3Uej0ebYnjmIWkia+E9VGi19KrhDCY67VgGb7OOQj0/+l
0kmGFC31Y7htnKf22l/vF6MRmRjg6zhDrK5aUwemqHMDvlb1dhkg61y8E2j4MLmL6PV5ZsamKjHQ
CSwjWpfo78T8976MiANm3N5nI6bMTMGU1fJ9xNrsG6xJWeMeGKgNROW5+rZtNpHM1rCcylh396H7
fZB93y56vLpIeiLWDArdRkn1X8fzQ/qwdWDqxs+HvBnHRf3pnHlzEiknuxjorpAoQHX1x1SIFWJb
m8wzAzae9/FqxRhxE0OHsaa52QNppKK+gyCidZhHmL9ua2nnBciUDRGHSsTecEkQxVJ5mSdHH2B9
IbR/pUWqUghMm88Rg57xsI6xOoH0uT8XDOtHnLMcS35MyX/8JCQiDrRCpD4TZah1bL59RjeepyCJ
O8RoxHJR8evwI5tge82uZkmyFjJLcn0wHKzrBWuEHiIw3thJl6yPoX4mRyt0AcPJcAKvF0szBluP
PvaL2eguDlJ35BlVVj9y8FHIs7j2tlWIbbEaedN1bwK+P3CSfmMfyV2q852wjr8fvAxPIEJ0uqxJ
POa7FV6BDdDVErpesAkH4kKVUNzzamGC4YVc0Fk90c618Lql0k18B1J4JEY3qFL8EnQYogYoE9Qd
iKmiQvL3+CIXQyLZpJrhHNEAFlw1/VtzRBRnXWTnWCUc6mESLNQrMWjth2LbbtCy3CNxKgCgs/yb
GJLxiPYQYC4xkU42bsi8693J1Z41qbzFGt2hAfht1AnPOJzFaZHDZrWicSuoD54WvEmVbs5ID/5B
Pt3DnISIxrMZJy+RKNWXx8ODXIbHisB0B/0yd4aa3Wgu7scoNF3glsmjCiVK31ld8LhFX6HwM6ht
azF4mBAtI1gyl1VvMOxvN34kvvQGviPogT9rWboDsP/CMpmPswnPuay6cJxrh+PC9hqxODhc/pH7
4p4z99tZc+I+uVOLXwypyGNCwnAxY2V81eik3e+gbLVsWL2j8VG207AiIMuC61RPmxjg+djtBAMv
ee8SrxEI4eYkXxNJZ+d4bSvldWGmDcouARxe8lZ9jT+OzIqIGNQHoTtvTFBwOBkR6s9vobJg4czN
4sHJ4kdGi3G04ralGKAqyTSjpDrT3fPAiwaLNIsyddfeNISukd1qJgq27hFIShwf8NOCX+iqbdZC
xVqv7fChzqbOIlqxmYSRHMaCqp0lAv01GkSmkmye9yMG74t4w5CJkwOrE2HjS4wSynOpTShsT+j0
eTNKP0bXSRDs8iU734f6qVXNq1qDeIkALYj8Zpuqij44aqgYgGrZIff7muVeYroGPcXCiNed7CNN
YOck6WZKFyC6U3n48bawmMgg4k0WMHukjcWuYnmDpMkCrF3EwH22ct3rItWJo/87mz0H+ikLfMu8
2iv7XSKdvNgnLA5sFuxEWE1bDEWWggYoImDfR+slFBwVmfLH7Hn3kVodAPMTAMMByjvg8DH65St5
HZ0Jto7U8ZH1ris7GuD+53NZ9xUrBIAvosVU47m6EMV/c1M415YGa68Q0p/snjLE8D09G1tmnVwr
rnpcRywp1bdyl+X6fpWEiy8Qty6P6A1u/v7v25eTjMxDDqzRth226qA2KTmWK1JMU3CBQmoFkHLZ
iByOgJIhCVGlNRTLhBf0u7VlV99wtsAmWOFSy+besT2xxyF3alelA3ZzLplon7udDgWU5hB1JFq5
jOpFkRa6KmejTuuo0qmquEo19EmVu9PMblp2LLJ0T4v7crPRn0+ipchuC0dsnMZuIZG+nXO8jXfO
ovz55t3Mw6BSilWjB0VxRzK0cdLOp3TmEt2QGlJCAbTXc14DFeDWXPea50eRfUyO8ed79jVYCG3y
mKP7rVpkGQADbc8iTKKjQ+AIrozpFkkHOJE/ebtvPYWK4P2UbzOEkSq7DTE/WyROpbpyfs5zrSkF
n5CDyf84RX33/Zr3f1gqB2/3QUkqt8auY8LMF0dAILp6VWy5HvZ1K14vdbWCfA6OkZtBZkdGpuON
1S0m6xLpP5eKP8qYcV25ZK0GV6ikPyBDZwXHwwaso6Bw7w6Ngr0gaTmbDNywREaCs/u0ZilrdS5A
vexifB77Mp9wM3Eb46OujUs/RalGlkE8975kNSgd2UpFbOO4/9wDr3BQ0Wm9nomec0FcWRmfOKCF
xVNaKC4gBrhzr3J9k4Q1UMOUm0Qe/O0Leas4UdlfyivOu0KHq3OzzlTHWzQLzMtkdeOkBrJn6BZF
VFIFLosU3bVhvfRInXEnJ8kd+FPCxdD8DHL+5+1A5rYLTSAzMzvmySRnzh118XJclmEUyYktiZUe
RMl4urrCKk781+H59xHqAZV+vYUX3AzjUggV5AJedmOkJWpXveSDG+fX4hyBcNEUHP0pnoVsaz2X
3M3+V3ozoQARpjrR/VBsAlRgMkG6nBkEG/bDZcrt5FDmxwzYxi/s5fkawi5ngbZxIKujF8vzuq89
MHoRcmjHyEOy+ktY9uPuXlgejcnwyn6GdLtXORHAQ/782oI17dmkzovvzrbFGCexibQix/PGvKlQ
SwWxilUjLnpr/mG0CCtn9jCmHGxzmGNFZYl2Y5XBBJwwXgAnaAyd8LpzFFqZ6Z9xxAGNp9wS5p8N
miF0itK9BvvOcQOdVzAAIGvA3w49+1LQIXL8qhWGu5cSdl6wq+J8tCah+olADhva+29oIyjL/SXz
7Ehjl8zFphOzFmvvcnAj2CdF588Zn7DbsHACWyflyknKEID+Bzc11v7kNsRhexp056hUX1+QS0MR
ZVKK3Q4GNF6F/u/XrQn1DVSywPWviAAyRn6m0mpKwqkmHmDU0dqHeXvWZTVfOsM5jGme6OPGp/VF
wmZFsLjJV6BkUfLSYYHBliFgnnxZeC9QkZ7RU+OxKyPyqc/hn008n3dt3hnmiShefcPlthB4XeeV
ES4jsHDA4SeX7usgzEF2dEAYI3nWg/nKAWuYCUb1XBQgfDPqOn2NFYXBD+lQyTQ688GZZlmmZ5Cv
PteDlQnkC6G2uCJkf4fxbFp2LMzFgHNczj7uwi4gGa8dSMDdcxAXbmwBI+KxMfOGg2ptabuAK/Ld
e4ToVvyrwxE84gSkmxNuEO4Q3SXjmD/xiiH57h/TVpvocAckrwKOBI335ECgtvSiFhrq3Aw46dxJ
JHgrGfOf5WelofbanuR/6XGNMpkMKs0s62PB406NiSU9+pDXLBjLA5ald8kEHvcHtrwyMIlpsyO4
6lACoQKXyKhx/iWaFBoceqgTCHJKLaf6bcuU6p/wfna+TcCoGNRpWgRdFlcYI6KX6MBIVWBpMU9o
3K9zBZUEYek4kQBp7odWiCVXAk3hWyf/tNxQxv1v7HPUuJHa5o25/nZW4KRuDvulDcY46QCTc9lX
oDl103PaA9qr8RU5FDm1HGK5DPfgq5tZgY9aipMpIUAM4tQFlR56w08ikRCkCmVo4lcBXmUKg5Gd
hlKJbMB/YJFfVGO3KhpEJex71FrYijdAqJlLcGnmslqAF2SDWX7tZ4osrsNHcNxcp0WT6BTjmeaD
WmTVjLsKH+wFIbbeR6Ye6d6RxU4vUqE6rQPby6dP4QK8J7dHx82bryyFTw5jMLvHg2hOsTgWjWcJ
oTLCqLdVn2dTEAIX08GbRiXRKIEGk3/+1C4bzZwOobnHnNQiyHz+UP//6gQLMqQUByxZLFBH85uI
SGVgIt3FmHRTw/vcAWJUvrOaTIpOQi6263cYiTibyrHhpm5LgU781N0J2GphSEY3lPfJHItdhmxl
06aor5kc/kjNQMWrqJeKV0maU9toJisWX11N2+KO30Vqpv+vzNGhoqFssleK8Fm1j/mlPaCmOxU7
f3KlXVXnfFimkhYUEG9VMV/xwMKzYal8g3ZfDh6OZS6Pb+eE0BTzCTLIEx3XLaq00W14yY8yeh1T
sjRlRzeGpzC1CWZd+SobDy+sMrHJmX25we7iw/emFVoXKL6RdWvrqV4lvcgaoDDZ4vTeIFohjo0x
kwhatMcSi99P9/7AYEiKrQaczwUTKhJR0uDJdmqJysrCdbsyjUxcBJx3o1zIeYsSwaNPBrXq68eB
GOOTtSDTrENpq2xmPT0foywFy3PKjTPxT+9VnlXNWCvjmSN7s2mQVQlJKxK8cSAnrjcH5Yxienl8
1TJCH9fCTeuBphv6KyWFxwKLqk3Zna3h5Faa3G6lo074P2HvgBnT/AbJvM5POTEBBCa/j3VuQZQU
yV676kJiGQJcqHFlLsDeItPn33rjTUWSj7+WvsHLKL0UA7gcLuCyO6AJ0uwUPdJkXLMjUTegnC7Y
9wGjU9rpV2DNUVyQeB5gGkiVMK6wsdIEMxsRo4XJrerJ6q4M2K25K9lXAS4yXZvVtJtwhp9f8pjA
CB2qAsd6NNCvTWVE9BpRyKaCAY9+7tIbTYtRh6o53iEvdTpTNqkNHp5O/BLfb/TXbMzOatRDgMk1
SU8MrTQni9MrB2BMl9OV7XEYLCgOvJsxN5oeexS9nWtZkhAGH9Gm+hnqI5XKk9oQ8kgexQSMTK4I
ZtnyNg75orqaX/JTWexOLqtSyfyUE/NbzDDR8C9dqsDxd/mnwvVVjorN9na2a0N0MwohGeLCv+50
lr4s2zFAvzRnLxaPPCm/x92NYxg4+hV+OAGAcX94R059w7IuJ33IAd+uGnWudvWpi30NYlWhwqFs
bdBxxA0trvGQb/e8kf/Lwu32gck3EICn+sBNjJGbsnaBAV/fwB02bLImBOUy7Ano5apJ1pIohd21
+lY6rbE6QhAtahnjoKk2Zu+pTCJyVhrDvGzg4iCsPxXwloBcaZYOS888NOe6DAGxBBom9l+9efxQ
oJp4Z4USTxgVVE5Ke+f4ZxGOBZjaWBO5FmKW164jWtMJKoibH0iFAn8xJuFlgfIC1FKPsZhj8FPk
UgImDOqEN9DRXp+y/LSYkKHvr6OkDJ6uifKYNI45Xv9Nkx2MqhU5ghKQ0JWMBm3zWZNyRUuIxPxG
9mc4IePiaX4TUgTQJEk9vWLOoFzJt4g3GnM/PCx9qI2RuXqJMgRzrQt7Fd2fr44gPxUdwvohTvxk
qMVgeowjPPhSs82JRGRVwqWoOtYcfBAZw/pctlgz3Sedtj613UmMkCK/kXx0Rzah6VbLBHprZBX7
xD1TrK7+vqDshTH5PUXoWiedAdgY4jxhGgB/kpTRa++vZKqnZNy9nQTkG5FYvaRvKLIXMqv4vZCW
GgJK6i4vUjhd7jg4slqKuTiD5iz0UBpVAvg7sbBS97v7I04cY2TMvrBn/RwO0KCKnrxfhjjYz7uP
PJcHS3NwweRvD/HacZj9XcpDp4McLcb0nKKG2lAPt6ma93WwjEfVZKp3eTrs6Co3chrXNzMvrjH0
iiRE/2VgaoMpT+jr+0zQtb5i0hGLp9m5sNZgMdYGIuTVlK9ET6nfRFaJwEXhW6d7SdiHIMy9hJIG
/Cpv4fzQvEiNePQHij4yHo5sDKhfRj2EaPTE7C+HCvXNfhpNX80FUP3iw4P/vjqbovCYijT7NW9n
jdRMrwWOBF2aeEOeZ2kbz/7BE0drzOsCJ3xCflIjTGxuah3xiAz9w6pHpdUuohh2ywlTNul8eHWb
7FxxwwdUFqKHbk7aU0wnjGflXe3q6XtZlbIVA1E5FoWlMfbo1MrumyN/xBpGBR0JErc43bYS5TMY
W1D5+R2kXrwYzwBslrQvVuxsK7V+cumqwmDrWc4/SNIYWQ0ZBxn8jg+kaM7GxZwkSXV9O7ZEep7L
Bo4E6bEecxTqhKQE0kkgxvmxYBB2YNDEsvT0Hm6SUKeEcBDHhuYgYNV/zolH//X87aKYkEL5E6Ol
xrJVOvNRJTcvqGCuj2plhpUJPyOPI72l8B1qQrH/xRtD7hoDYfoQer8IBXEjDa9NmH32VpczYfov
rN8Aw0Z9+d8T8Ghk/A4kU+T/p1Oz8OWFUBviLj1m/WAij5uFJVWn0wSXI99YDrdd4KoC0B8v9gns
13ObDE1QxS0KVNKcOSlcWtBSCLpOD1w7gXqh8/9eQtiyUshlrtXq6/JlGdOAvhbw/MppU2i5UuOc
HkY8z5Qdevu5aasj+fKavYOWku2pI9er3sxePJiWMn7J0DkASeKyWHSsbEJZAhJZgdJ9H04iT28J
r0vLWahbFzbxoybY9x9CXZl48BLMDJna0/IzbMrtZYaoSCLPA4U5lN6Bt2ceSWzNN2MMdV2Km/LN
TpQaiTWP14Ps1dogE4RfIST8rpswrDArF8yAfQdgBcXs/dwO5hUm5od2vWx5hpBySie2BzE+IIg6
KDTbPlAbCwW86GJ4uU1O+2jLsPW68kS7dQJYNvkBc6ireR6RcEwwFYoTjolilPOBo7GufbqnfNRR
lrWeKXtD7FwKDda6yNfzQ/1UicrZV+0EWn8yp+psWKgprwYngQCoyRDaXnR9Ze6N96Z99Q6tDDAh
mauaSl/us4DmYG+xrY83cPpSrRyA7AyYpl7P3i8R5t7NSJ9gahBHLonB2WElXST/C8a5yAXfl/r3
6JXvkVCdC2baYE7dez+RXl3zqrY6uLPMR8kUoj0xm9gQF8/PXj6ylwUhIH97Lmb1BzeqjlN92wCp
Etgq9kKS1VCTHIO+EYIW8NL5mM3hhbEaroFphhUPeKUq6Qh3bNLHkf3/y5m5Et1oyptb/tSSKMLE
kiKW8SKioQw9ac+PGbIKhU0wVJ6iocXJ0qA+yuUbyo8Al7UTeZf0LQC7d5KiXXQIO3Leqy/C7E7F
8favnO6C5Z2DRg3p297HIeto5Omvq7VSGTz+7WgodWTzOxfjmPLocVwApo/wOwptL26hs5FopXdx
qmX+Y0YCPgaZj37JJiwSFOZ5IV17j27qOU1y9LWQvup/m/DhTr+tSfLvPebJKrgOngYgSPC4eFCv
n+cfasC4VNl4msWMbGWRqD+vpW7sa9KDWBzkcM2HNAp1BFn76QFQc0I8Ke3pRXTx7h31Rq5eX+sI
Zl7oA0mkEMNkN2S5APhj9s+a10wo8mGxkCp56ovc+syb6TxzYosNOmq3cA0n8Es/k8frdE6rJSWN
9r7oFdbzCidDYPOMJW5ymQ/ju+fSkxTf8LtHC5rJ6vQ4Xo4U+pE/6ukKIXGq3lJPKlmKCbFNv2XU
WP+Aj8NGsAwAb2pPje0ot6idiWZAadpqKgJqtvLxV6lvZk5WFduZQtBZYwQoJiRd4ZLvET+hy+WM
sn/xoNNhsP2Rd8z90XlqJI4N1HuNlfe1NUf9g/OFWq0msFQGX4sa7uQShdZTubzP1g4O1AMhl2hI
ktY6K+HnejBsk2rG3UpLY9e/j03LLLYK34WB1+skZfi+cyicrJsZArUx2f+M506+satvuTapGiUM
vLbNc3kPeNpu/3YmUlqSmuj4T6r8Ln4ybf0jOg+s0oZIJc9aDw6o3+faQxKpBXKtkqsrDicWguMb
s0tr2olejNiOdVJK2eL36Ne5xlA1XKmrYdgKijN/WBk2P0JoDZvqDaPpubmUvb4Bz/u+5TrZwPBs
oV84DIDPJMMAJHXutkz3STsdMAZDCuLSCkWtUT8Mt4oamJJnLT9S6qDyKjzgzCtXKaJwICflsYhP
xWaSGR8EjW7VqXS5a743Lzo5jgtnQ9T6Pd0I98dAbVmdBnGePNydFAwBWIym1NXxnIxMqT3bUqDY
Zk5pXg4H6SuY+zLxjYWaTeyjbicaKK+afYOzMvHFmZE/ZeCImxsZaJKUytrdeUIG0SAR0egjvLDe
sjcj3Lo26FfOhWSZQ5isyxaQ60fZGnf7oWV56SmhB2f2Kn+iLmWc8DCcP9Z005LauQXwnlPpk9vX
ExhPKeu0Ged+GZA+EY1KUkTu+OZdsmxPkeC2lq7YiWjBkzPFWvucKqe+HbLrb0ggI/K/h5cpt6eF
cluv2Z6Va2qOJzhMu/L5gFVh2gTIu879Khh7GL6C1fqR5uTJVJ6csyn/8LEDHujonJSPotKviRSk
es0NoN+jkrAb/vqq2rTXR7qiiVIejzNIBTZ0Xv3Uk7jtd9c4XvUdzehzg704KzGA5Hyw3Bsr2SJP
yYl2NKC3hE9KLr6+ql/3qocKz9a1MRwOvzTqRDwOML43EkItB0xwScABZi9rTl9W3ZbQkNAIOClW
u7wdElv5Q93Wur56EgqlUCc/O1xP1gEKw3fIXp2NenQ+BUMylFlcHLtI7bSrEvDTmTqYB0mrwf3b
IrFZk+k5BOv4KuI6Uye0p9JQrlgR3nh0V5t8cTdhjBvTug15h8xen6lyDiSGOebLMPi6moI9KUbv
kuPtrN6r7k9wAT7/0lwu2dW+QtRyXT/r5NqFgAcTqqYiS9y1kutqQzpp+624bMCm0zhNMdDc2qlD
15RGZEYB3yZW2be4Vi5uW7XVBNaGCNuzP+Jm8g7Ari6Lfquc7X40IcR+ZWhk7VnfsTafnuvx7IoL
CuuHEx8oURdC9sJiBqWTVzxA/ue6baMQxqdPfPN1FtaPtC7THNJr8pItncfMY/KZMOd1IyR0nLB7
isCI+ycyUogjHLJxPcGuL3ViVMOW5HWyGZzYEck21umEbf6CDGIq22vEmU66VTJ/8AfxP+TaYDDu
f7w/r4Ofa4lrKMz6KPUwLC2kWoAr3eCOk8+ipJaKyUukvJSUwiQrUqcRYCUK0/bqIThsg7fugTlX
6GgwtVHNIOPa8HMj7xGxwmrYAlZFCe1EQSwm/eIGZ1S+cH9GI13gNmFjxX9+CZfkaLiXcmIJFKr3
MFMc3LMu7LXXd/AjnQwd7pqpExBBQk4HjVgw5kgb1Lz508wGmgGdpCBpiKEQxrhrVl9ko9KwjGUI
UJyI47ChJxwhh341QRItxHdgeoyBdPAa8dmXstybbYlOfd8gLk/qguTQHqqZwtWKYSX9OlYnR6yy
bEGup+1RumoyRV0YQSGwK16uC6Q1Tjft++u01db4zOXuT9kGkgINJ/rgkUbwT7aFnEl+37Ew+V8T
PfifSVqiP5FdjjXjpWkvUsROA+7SY//tAhXOIsxmWz4BYx1jItSXAjgDFM+0tF2Md1xTqhx65WBx
k3cP5GMg6ZZSG1gvbcJKrKkz51GjE4DkrQUIrH3O+uh0FtPzMzUa1/L46IwDHDgTps9jBxDDdITl
UQ6e0UBiHDKbikf0WYkdoPSkcTMuXFZmOByMXIL7JcaBhJTU22BawBwfD4UNsHiyS/M4svoa+LJ5
cNXI8EGfIZHLMBKzSxa2imqr4NeRkAlcpp+O+CSwmPpHg4KPC2o3iSU9LNKm48q8UwvL+62TZqIV
lmSSV9LOGgzF6XZYRQkiJ+bpO4zBic+MRTRgS8URXGIhe+eyPnQc2zqVEGJOMO5EQ8sZH3KoAnbO
yR2LTpaJzg+YASp4BBPzbZ9zZb4KDRc+Ts8lnbVMD7Yy5oOPH70mzuLogviVPRVzP6zFBCGA5RNP
2W0mUASK8C5Tw/LBRJn/a4pO3jTbGzkBID0zDADvyORpBVF2hQ5i2pvfCzT/JhCkwUGDXCk8d5Qx
cFp7lB0HDv8jA9gJeJYYojIiWqObGXwCVgAXxY1oP5RHWXR117B2l4GyWg0JpU0NjDypgpBwEwHu
aHQ6tbetwELVfZbiOnmILOYqKtwg7UFOt31BK8PZygkW3JxkuUKZCaPNoDX2AYzuBREPoWMi+fGF
KucbTuY8yKXuZ+JpCWrIM6e0KIJXQxYwc7vNBGm/W5EZ6ho6DcuOSij0JINthSeJh3/BLF030AqQ
zE+pPYkwR5uVu4CiZQ6S09Kzn4vIrxzWoT5Z31LCr5OBl2+P5jEH2Bzpz47CI//qPO7MddlEuzlU
v+o1T4wIi6bn+lsctgonuvcNzZ643s9j3g2Kktwp3Gm+ZqDUCjJ3zRD1Ctcfwrv/oLCkaM2KPihZ
muAWBsWqtPEFdO3UTiwaIoK/co+D9JQxc0pETNnMD1tj/5SvPuGfqGW/xPzsuCxXs3CyjmmuILwJ
6bmuDhUdNxb5XmgBVCT1tufZppjWSct8cZpE7ymjjYooCqSun82+2db1JL2IxHYJxlQg9OjkWR8o
7HZoiyTAeqKG9ta7TdUlgffw7OKhInQqexZ7QTayy9LpTqgDxq7aDeAWP7ATk/FueCNs4PDJVUCA
zEVYk4496bQ1+xFNqB2ogoxwlHG+C97uHSn70z9EIntOv84uvM752R7equczpIEc4UGSlQ4+S0Ly
8/PBxNETNpWBOtStM05cxKFfd0CQeDxD1U0pk7GHS/1VwVTRxxVbI5EKF6sIdRvITUd/Kr+xLoJK
6vTWgIM3woyq92zHx9UxEMYJ2A5xQDv0whFiEzdbafsXCt4whe5k/0VskMyunw5Tyi9tTef2x3qb
PmuyxyzoQ/B8F3UjTGYiaeLUSg8V2vUTwfZ30sOJ7zkEILFHRvWr/ZlBWSZsOIqIQe7ES5s25qN0
J5JaTssWPvcxQdgIGqkK8RBUe8yrQ8J7DzMyEnD1V+kqNlLXbZozjOuwy0hlWytAhH6ZQnJ8FxBz
/Olt3xZs9xYKq3Ax/otnvGla+69lM6gjs5sBjnsfuOI7ukXExGn+P7iy+hKn10u1GV5Uow2cSS9C
N7d7/h8zoa2DG4sJ+vFxsCSoJqaSBsphqvOIaRTgYsJP5gSRb+ch6/P6TL+Z18hg+IbR2O7K+E42
aUQay5MyIEpavSelkzFxtL+CxmjTl2/DCVduRm48Gm3ZVD8F3Av8cnRlYYTDm+d0A3+VJ2OwyTUZ
mI//h0Y8niu5+q+Uf5NO4y3QEWqZGj+ip/xdZQs9SozlBN0gzZ9X0rlY7WT8gMFlTcKCzg3vZim+
HMGYuShyROk3nBIu7/iO/TddHYF6WaP6+88bSWrMvFAtNU8sdz7lFJ+3Gt7GbgnFN9IoyxFZ3ubl
EEdJ8KSQ+vUBtjAq2MFvbGUNQaE2ARNUdCWyoheC633X+HfqkpY2wfEhUWSLaxWERCMBXnyQG1zc
E/lyFQg//6JEaC7FWskyl9Y1dITH3AeIqqystBnwcyJ4Gwh670XvBbrWn2oAWaLDJGGy5HoYFPEg
z3xPo4bbJktm+LHmHVZmFEsd9soA1OecWg7ai+wc2xpOIg9KyY+bhoXRYzlYTkAJh1mjTRwaMexJ
SD0WQLQPeWhzGhr/cUiWzObolJKTEmDJMRM0QDFw7rUJJQukAK7Vn7HiX0pM0JKRIkIUwEiekDBc
oWrQjmlRmz3F0XsK3qlXrO9uYyMcM/TM1CdlFRffHfeGpIlShnL0EcKJK/lSlJ/p16quXvkvP2xz
5UoROz/t03npPbZonY+XznhWG952TE+amqEg/fLHZgn2UH5KI7PPbG+E4KXYys++9/HPwv9IE+0E
fJwn+AnIz5TH0kUpQXFrcmYf0RrnbPvcCYnGO5Hh94vbomxmArWV6RRYXHIozOTaAetcK7N1yL7L
aYKR2t4ZgoLSs3RRPMEdy+SWUauwduZF/D0Qor42lY45sNpau2y5LkIlnafrvkXVHPqIAxa6bXkY
kzALHdsdUlYIyL/FMY96/aL1tnAPykoMbOqCHOLtSQ66xFlS0esGmWDyB8mma1jZkgO0NCRupI1l
2xcDIL3L53GVbNNtVzpiIP4YIdb6daHDxxs0b8luzO5srONh3Wr4lzE3B2Rd0JY8wJGIz77TZ8kS
/4fxWlflYC7fBcA7FQ3rNFySxOF9ZKkcfhxOtG3HSadbi9zZfwY3f0EwsC+wbAnG6T7Xa0nEUthH
GfcCOj77D8nuwJW/FFZ6iDgbjAFRkhpFTYHaYLxNeUbMBs2SO6iE9MGpAmq1FZx5XiRO1+H9uWoX
4pszbeYk7pBEZeySOZlJV6CAX0hx0wpRrvzLZ5JeN0z9CiCql1Pp0VBgZUVMS81bb2AatiXId/gk
ktvQwcmUIaoXYZA9oK32iW4SDP3V32EcKXGG9sLRCHBYyp6cqwcebSgOxMBTgjFlYZMx08Ns85dA
hYPdJUdvDz8kk1ly44KY1ECrq8H1TdnG54JiglPkvGofaOUpxzK9ai30fpOJKjSABZf3AVjuyI2K
d7AQGUu0FSMcQldDmxGHTtWRvz4jyGxhpG3o8oUoldMaPe1f5JXh8m7sKwtP8AL2tWh9rnkmV4an
gAVv5k9Or+3jtLj34rC/8EH38o1RBD9yD3zB4zQj5A+eNXzqbN71xtPV5Ka8Y5ZcPSVmR8wzU1iT
+qzfzy6UcJJPSzU7T0JLAPZjTtpB250Ok4EtZ8neRRg5uRPXr2WxurO1Y7ZL/O49CRSVPn1XdJTh
Mmk12ivwo6AEzFCQ0Q6O+L812X5xKs2ILleJKLNsX06uAVsdmIB+YIkLxapcIzrFEiMyrnf4/K3F
PN5aS0/LQWsrEDIROO6zk//CzcYEF7YYKpQLsb6UgXrGXcgxPgzm4OOK6NXFOAX6ML4Qa0/49DLo
FHVcExeRDKYSpViY7EA0oZVYX93yPgEnm13MKDOjmFg4YmAzfgCA/d3GC3GuIsVLpuVRSpUmEsYf
wPetbvGJ6iZHocIbFTG0QHI80BUw9sDOzuRrTuxPX70f0bEm70SduAhJ/AmW0HTjRj3S4y5uP5UB
S0ggMmuNO6r8zfuLc90g7IfAfyw34vLagZ0yDIWSkygPWeGtKnP/Yx9ULpwEwIcuOfmONaJcJimk
01rDYT+Pg7ve+KuWSFVupHqz1jAjmfVmyXCtncBFdZayovfWuXVYC1BdeHRCrG0bd5WAl4MnYriA
9IHY7WZpar5dLBnjqP6FjPs8I+DvE8RfnYVro0/0Y0xSIGen7AeNW1KhWjB0TGK7ZIXx5Q7MyEC5
+TtRSyX/JhaThCEYe2+xl3oHYjkV2uoOAyTWNEbg1ECJ18XRnc6fIkd1XTYN/XoowUgs/9iX3md8
a6zsJGaxQSpWZaFI2Y4hgoFh8L4QckfLEEJTrrRxEKNboFvF9sMCfK9Fb3RsAkOG/rhkPlB0jQlp
pFegMe0ENYSak5yvJ3InlUIAdkRP7aYM3lofUrrdcSgHbzib5UGfSQwb4ZL5eiEIO3E/p4x75exJ
SMV3VG43Bnf0iNyZKEzLmkDAIRQcJyfx3AHbAq49/WBRhQa4KWC01eumbaah7b7d886ZYYBIlTbQ
X3I0vz+X7Xax32Bk49HihSFxn2V/IS5terkYGKzaQFB13L906DuZjBYEHT0ZYvrZqSEDFwWJCmR/
c2uSRNg88/4PM/O6wqhGcB+8RUmBbhoEmPLvtduuc5MuwpmLI6mghING61onEZtwhx13VVqlnzGl
YNCQh/tX+PFrsVE8tSSkV4bC82Dct2RiaeWJEyatqnJEY7JzUEaeIoz/wie9PN8L+uzN22PNcSFb
6u9uz1G8GbQ5C7UM10zK873F5OF02V48fksbY5thH6W9C9hR2nHPM+tjSzO1jLKDp3u/qMEV868F
au+bEqD6qDkEkRs7X+8mraezb4icBauULqta5rzuYuyn+8cAGU6m+ZVhnVy8RFJmOnVZ37FA7xRG
e35SV0yxulp8rNDjvQIj6OajJi4rMmjZeY10HfgnJgfdt/kF+b7HG1Vqzk+qGQprDUlSfPCTT4Hr
USRaXzBsAbhIJUdX2m31PdwvdOyReczz1vJCCOGfLcZpia5wkhJk9+ifQ1uudUN8MZznsBE83I+B
ErWdJ5dx/ktsB+soMnojCBizgSZGgrrcZifowYjFQSB9MFyB4aV3o2cqtnN2eF0nL5RKxwXHR+kj
JtdA5QyRP//wZuRrQj81YSIE9GeXdNn7+uGYX1fDJCS4A6E1FOctF0Z2OYtbmlejYPNpoJi4Fs2d
tN5dOqqFnqS0pBnk9nZWsm7yjr2Y7ygGskEPcnFt0atsJPkyiRyYpXo4gf7lwjEsic3YZLKuRTJE
wfAf9H8jfC0ENFdGpqmMEw+Vy1VRfUlwt+04DHYNk9mqzY6GFujE+amJTX2Xmf28B34ZiiSdHvc3
R3my4QM4tKaColvffbVY/Id8JAhxSKvsDO7Za5dpS/TlaV+0pwWa8xedXIUl1icKZjW7tZmjNRLF
HhItnRjgMVlmvQMYC7tGq65677AZgiQQGhQi4Ea5zG5mXXGz1Q/KqPTYBjdR6wEia66CG+TV4uyj
V0ZVvBuF1De7Vhk+2+uFk4z2yGjATcYA+IjDc2j96P2C5R+ZcXy+ssI87O3NuQ6/9Bp8PDzAUWhf
C9VKqKWMmDGUE5D3PrLd/J5+3ceHk4D7VZOfE5QCovKqlZp5NaTyo1hzAFulx5gzftrUYPVeYvnS
Q6uNZyhj6yX415xclqqb4IBBJjHfgV2Jx59saXCrymDn1M2s37RsAmhSzYjDg6FHH9bOZdXp4C/2
zLoLSWAA8QuxVhHKV6dX6vIaeKiAYZ4+Q3ZyA4wdN9Lg3IjWo9iFGLwLDYbGDypcP3v6whLcoBrI
dPmeXF9wEJfO+MwIw20SiWNixg1d1jzHzXs7Kg25NYm0mVgRNheVojJ8UIGnCrySEaWY4Cl+q1kK
V+YRzIWwxU6tS9ixpLUUOnVjpXqc2uQeHLzCCQpa2FVPjjAqZGm4Lx1FL2mk1H7fl70LJkcrnnn/
FsvczM4crbad591qm1vsh2XASp3hhju+rnH4Bky63OEVrYU8Ke9eUD4nIhow4FXSpbE/I7roR97S
5ydP2XTPeJej13imk+P61o2ycmCxNPhX8B5VVim/NWnw+J7KMhFgVCi5ZjLWepDO9e/yjS81eMo7
4hV0skRSYHMc+jYyCCceROlLpqzudf9bONYFhrAlKsU0TeS8hkLIPyR2Xi2NW/zXOR6KonEhEsXW
FigFMcKb2Z5Ie3SFSkCODTvMDBkDklk/VON9R4yDUlGtLtyUHEyPsLhT9Nk+oo3LEYeB7iiaaiKg
vF8qmlMzErsBGYp+Rl8epWbx3jBYjuz0X2QGknTbwcSUZ5cLHieuUcSbTYg9tShpFstVt+1cJHUl
Y58TcTknPfJ4QRxlSvN6oxw2/NdQTCTnf/k52IUglI2d2Ix/UpIpLHlUSNcTDA/HR8m/YwwXIdfm
kqebYWiEdZd6Yij87qIjMc9jlOCUHcyE1Lt38nzHW4b6VNVu3VhROeZzuhPNhRk6U5VCC4dMM41v
6W7x7L6Hi2R98/nuCdlJHt95IHtd2FZ9YS1KNF6C5grPrvFAZgyiBiX8QjbSmftkzd5whSyfb6Cw
a2GAWc/gm0WfwllJTowk6MeAsxCWePZPMJN/IpNYekJyumSqrou5aJizrdOy+ygSHSnnp1LE2INu
kXGy8kygnoXCWJePjLCGIcXsLobtwXVhyQOSdPd8o1B16Dp03L3xo0X0a7jcmam2atNGhB5q20bw
o83QxbSWCEqoMcUoXl6Mj1r0kk1kb4knMmf2KlabF4eUo2YReEj1CCBZ6aTcX+wsxwJId+17l0B5
EZ/Tm4pf0290XGYt5nbPLUM6wWhmk9hBAaOupEVaj/11RBEhCa/ueZLsa4pE2S39PHhRbpmNo6gO
XUCHX/Ch3vKWGVWuViLxiqnF9+Xt6JHuMMlprFi2ii/C4puZ2X1niZeSccZMsn9DN9rQIPiLd0b8
g9lsKeMHA6j7BMnRB+OLiqyvWABQ/l/kDiYv5oD2MxOKWtphEkdAWD5UaKXI5po8yRPrcsbYQr6c
NhXhPR2U27hpWx8/zovfj7I/B4MTFI3SmiczdKajONEWioGMl9bPoFRvEHzZQ1dtkshlMCFgPbSp
YwuTznZs0FsK7cp8PLBpMqQxR7yd2jrobO9t/Q6jpYbHwTWsAmpHIoPXM3RzQ4Me5HZH+5pkJrQf
H+VNizUwB0Hz4YmHe8DBwWAaFQvjF0W/tni9bJXtS+za0aCibmhG075diOnqRbfNKkMy6pMA65fx
hTO4rj8bMlzXCcUuzqeFmKjkP66k6boRnW9XJE5gxbLKfitbHy1mnpthPUGYh5ebMzn9WvgyxSut
hEJkTa5/fL9VZMPi1/VtxzFc/sXwaaAR3Ufll9YXE/Wdpkw68tWIRpdulU9VlF0K5wt+C5OQ/sWG
BRoxgQoqgkjCt9WSLEp9j3IuXlK0IRZ3AXX3RDQOAtSh/mH1vr902Hoo3wBq8A8r92wRfODHagIA
P9qPDy00HTZuN9MJgWji0EvkG1GjnMWpLxLt559L1ht0aehIf9BXUR/vf89AZ8973JPp9+Lni1m/
lKUny+gUnjDtkxvjQHHBJPDrFly6fDIV68cMLxMAuY5+7C1eqYO2qaATSxXcrOcwhWP5C8MylcBy
r67rIvhP/+JgNPNGuohai3xPsPUShbMQUhn4H3yLlu3OEqmiHRyRJfL/A4ySJrAafDwgZr9kXPoh
EzSsUEGnxKEqr0Ki0dyGHa4CnxgvAFXh/Re2U6mkQFejp+jCpsMCkafVjvr5axHVsUuUYxh37Qii
4i5VF5XJwmIG7QaZam75Vzb2Zt0Qtuvn2rch/dF9KrGF/VxZKGJQWlyo9ESsgB1UQncZ6Vw3Vetb
yAWo2VagFFX3F2G+rd3kXr86XE+DixO11THp4HmX0Ayg1gX6qdg13LWsirHxEuMCeE13MJ7JOc6U
mTibOnf3Ns/rUlXTwL4tFFj8ehRAQNWEVOvMtxmWJx4em8wqgVrd08eJ343yWDK8g14dNhnpSXj7
jwH5/8QEjem+f5eQfXzCSUsBP1UKZmKKZVetEDCy7bcYeMmNK9sE1sUh5mDd9RbA5JMTbBIDNiai
jhwa5hb3OuzPmEIFU6emQEHPFia0wR7vc625nJTqJ8eazT8p3dKcv/pc6zclE/uFeWyGMXGTQFH9
yBVXFu3Ke3nY6O+thMgLwIZh3Rg8is5byD5vXzFAV0ZCaHMFDo5ZmBVBLkPtYuMxbYwpDg5SqSZT
s2ctHFIL+SVqJyxyT29f/RYXdsHhwC+xjcRnHGwePF5wTh1rHDR5xz33l2T29fwILmGlWE1Eyf4v
ryeMVZHbneOO+ZbTHRSQl9IOxZB6y/uMn6tuB9I1ItACJOL2lMtKowk8k82S4Zrq9BTDXHNkj1EM
9nRsO5yjPavDpli8NNk33buNV3XQTTe6d5W004VYJvLZfYG4hdxwNDhefekgNH+h/aMJNtuuBtkV
wRypMlomagQgw1qDre7VB1iVVqNHMGbFMv2J1b2utqWaGozF+lhbSM4nyTbVhDJr1DDm87q+STS8
xe7e0CiROzX2LCnQk7Al2N7Bnfz2RyxQwVvNsuJSzcfB8Bxt5KGXlGirbuW/JZtD2X0VoiSI2K2Y
L+C+zWzeyEpnLbtk2fz8P0S2yRsi8mprK6YFq5rN9ye4NdKAec0lkKGRDxGXo3rgzP/M0fM5Wp4Y
7giylfOMH3bRIFL2KOWuWPGAfiJSc4TI1rqsxo1cmT49xkyY0bveaIm4Ca3nqIHlE6YfeBBNv0f3
+twQzwYQHqgU/Reb7aAQODGwzTDM28tGZ8ZYTSJpKok+12NMtG1nOezqN4hTApMiu2fRo3HnjIbd
fai/JuZFLcQ3W0hS6pvluEfvZy9+RWPdhbldA9yaUey27Zl5pCVV5n+NKeory8TCdBXDsF3St4/K
039gWBSnrA4ZErURu32U1RKAuMttJi6hfkhEyaRWC8oX29yc7OMDEc09A0cx2sEi90I2lYKk5leZ
lG7JGM7X/mbF7Vp/jh6ahMwFT2zFyVPpisK6t/O7WWJa2tx0jCB1YO3Ok66om2Dlmv32KBc42vqF
cqaCA8khVrscR9R4fQJeON5zAIhaY06t0KAvgXYAiAshgjC+YI0P8b286ViTmekdoLQNDpjo9FgT
UHsI1QzKlHT3qYApIca4REcnGdJ6Un2RrYBazJ5w8J77LLS8zkEVJ89HeauYdlwSHfHytt9UN3Gf
sSxohR0pZUGH8+M4Acjh9kw8S8QCVfq3154GzeU/QPyaCGOVsn7I/ke3xJcm1builgiH61vqi3ax
78afOgAppg2yYcnYKP3r6lH9mLSUgQ0wYIX2UjP0qN8YS8Y7Exp1VoL7MS3X/YPDFrFb7WsIrv5n
aRYLn9DJHVDTzbZGR7KIBy88tID0P0mb5aZDqSzwq1yhzWNwbZbKbrCb3teE7cPtx4GXTBuIC8XC
C9Bk8oNmV3iBJj78HMk8oah1dXaxCUAEpImxBM7eGczhFwEh0OZnk1N+acgxdnn0HyzFHz8dcsrZ
lj0Er8K6o06D5szrZtuvb3edC6nO0U/bok8MEwwwdVm7Tyni6pIzyfX109Ad8E4WBZ78ijZn7n3N
wjG8jdlrqSOfjK7yQLHOGxi7gw6lwpSugxdp7T+6mz8wPnrlPe0dMjhFe6RzJKybGAQZa+jjcC3j
kN9G5ePlg890Y5YqXNBBOoE40gfz1ckAafDmAGEKIzQ3QUBmKMmlqfJn80K3efaGRaRb2QbX/b8O
XsiNdCQlIYZIOuTjta+1gvZgeOucODbgoPk+zLN/De6S9+mUn32oGCRZmdejouqOeKZlDZpcLlMv
rc0GyNm89MgraBAGb8KPKI62XpxbR9YI3iIb4p2KmAh3NWkeyZPJOrWTTUosGNFeCKkNkZsI5ZMj
OhT0tcf5idOJzMBDVPmV6DrERG65oEz1MiGCjCpkpC9JdlGP358R41hkPZf6bZOu349GGgxQBtRv
ZYo+ML603fvWLkTwY6LlMVPtrpKsE7qDKXSiJBNlpiff1J+SPpDpiIvABEiykDJUQFuOUsTP9DgS
iQCO244WHuG1M1+lvqyaXaRcqHQIvFOHzLja8hgdJcf8mxtChq/iF6CEPEOwZMPkZVphBXiWcKLi
hQ3+wVgRW0RDZeJgexgzNDC9DsGREV3uYeUUb//WCtJB6x25B6ZsN9moUFpV9xe+kRpx4172vJ7H
MG9ViLiETXObN2prJt6p3nn6w+TalNVOwp433OSHgZQMxobUyIoeT7HMZAoGi01OG+2cmnnfBdZx
y5oREhoy+QFdIBz999gQiUSgtpcPG+uAlSQVZKkXwa0qwlceBoqnYO9iDGanSmyBmu/kQYM+WwPW
BtY4tD3lUK8f++aSVeU3d8i2nQmqQCQI2eI4CkKw8Js5yOcJTTvEsAxlh4VFnOPRkVh3e/2UWn5H
0D6jIfpG0JqND1l1mry/qHcNWNNtpBCyGI0RV0gn0ZPtmeR2Et268BW/fWdvVoe1DhlTf11rvTEX
a/+r3lP5CMq/4UYUQENFhgXB69ufPm6VP9mzXVYEgie7xFO2AlH9W1fdZjSUYplAHsgxUzJJiCuY
ALbdvPYItnAu0GTt1qsyczlmwU2v49TO/DJnSbE/87nzBx0z54HdndkkfwWOfETFzbDIvgkZ2Q3e
d2Swev+dNY0ZWeh11xSw0HQjrFyhgv4EHby/Tft49D3pIKIzhb2PeKhm9rCGbh3hsR/SCZ5s9Yam
3+5m7+cYJmS2LWiP5Me8DEA6abs5bdfATdDfGBOgjOWnhpuQRYEb0ZZxPJKkyun9NWHX4XPMJT7t
7sDfB0nqwQZPjnDSug9+fRsGc5dt+mM3ZJBylKwbdHPqZQNYUKVmkFeX4Yy5ygJ4OLFQv9RcKiHL
uAUNqnNgQ5vQJ2KOSgfjKY0PHf2Lq8XXxh7+Q5iAkpSBOhQ6VMTW7PPiFF8rRKdBHImNtrFHy6K0
HkGd0m4u7lwUk793KhdvZ2sW7xSqW09mwo5RgmUm+Pys2EpaQ0L0s9h0ameb/hyo7J+xZKXJSnjr
7f8gcpyFRcjjwNCzqAuL9nbEIjAfSnsnnsRNWcsLR55+a+6vuP0/HZuFm5x9KNAl0Net5q1urkMd
lEWUHLF5nZoiwRxcRdtQh0c5Bsql0Hj6yBxM3lrpY8fhODQb3hVFQIgr84WSM++PS476zOVyX8MZ
vttFrmGRsL49/OtlfXcDItEemOXmWdQsLzt7jR003WBPOZ+n5kso052ba47etKLU4Snb6RD1QdFq
4ADMduqMKAyX11r3WTZgDeJMU4FLpz5PAQQmqkdx2VwFgRTdDfhuwPkyxhS2/xokf1fwf5YYlCBX
9wVZfad5xqFQW+/ttPUib1+PbHke9Emm6ODSHV8nxDxLZKQDYpOR1f/RUhjdsWlZ9EQgM7miT3j7
mBGD23BXzLA90vGw4avtNCsY56jSJuGXZRysqNsoHRr4/xm8vrYcS8dHjq4Y/Q74tXNFBLer51Od
qaJECH6hvLJYyg3rVpF0FM7y+AfzofY37ba9bPo7cym30E5vrl/VciZbRWOAS3zdLVTAXBRf37l4
vl4KR5+E/MJXSmZAOcTOll72g6aoc28Dpe9RlUzjfp7lDBnLzT0U802bDiVRiTjGYHzoTbU40TVa
59+2C1r0Y0gCpFlJcvAWvbxep7ByOAef1pXmhUBBZ2jXVTovL+h+pYBQh8m/rYJfEkqGoDhvNgsV
XogsOu+WtEP1J6WDXfXVWzn0UwA0sH7JD1FXAqsuQInX994JXyb8nquGRoU29TBZ3wU1fLYhMc39
q+1D/2V22tCxaLfhA6paHaoczvpDXVMtjPWYd/5fs466Jgp7ZM9d3kB8A5aivfD0SfrsTHhdnM0F
AtgwBeOpiWmZuuznjDAX/87GK0Qlit/HFRpmLzLxSbR+qF3GybGsGNEvAiI8hMzDgPN3dPrCPJ2F
vSijAYRRLGCp2eGVf93H+Ewo3aGWrCfqRg5nFtVUH5nQ7vDKN7FmyLb7IWhPqmSiQhzmHaBuWMSQ
Dq2ao/MZiHXn4kSmHX9X1EiuhLDRFbyro18grC9zqX1kRjcOg+LFf9LdxXD9jkMeKcWVSTs8TZzA
QUMzET0uqsnZcDD659gsuyv1JuQPOQHraovJy53z8onSqHkpUWIavbqYEQvG65/X8i8IQx1WRMaU
I6SH2HtZk/PHb2smjjt48IuPNySIvdHD4axHNR71M0HMBviWDbMxNT8dRlSPJgutx5NJLHZfDmIn
WBF+HbuMoBcn6FR8joVIFvlEEz4xHQn59q/jJxTdoWf3nVojn9UbtvjiZCgptDDX5XxVJFB6svIS
glnwtAXp501RiF4LEZihMx2XGuT6tGlIq0E80mgbYdleZjBOHIDzsJhz0OVxaIiwtZtsGXUDZZMh
2bbDp4TYV2zD9/XBp6gvtdlOTlXv6itQZ1o0FAKvswh+Yv4TG0Gi9FqlVGpDAcE2KO7EihzF0vP7
V4D/6AY6yTJOeYLMv9HnewOQZLzLg9Im0zjiAVygkfBJTZln76EN66SfW6yXeTIkHTAO3WtC7LB8
u/IxR5EYCZFg8luCHn+TItEFlhKDVdKH9DtGc2v9LzKV8dtndwaOWNncM38WaSUZJUvCz1SucDcs
siAysRtr9+oIgmiDadhnwG7jFSfBJ2MC+ghkJ5vpJETW1CrKg0rENc4ec7Px9sPThAn4iVhlSXDp
V5i1Toq/LP46B9oVWhF7cCOUYlmXlsinnSjYIprPtvF4Pln4hJiNq0tv3Y4bfCSwbeV1JOjQtPVV
ML2fdykaNGTL0lfmXpuNUlfExwE5pz7UP1db90/za3jZ/mLj/9MpgDgKK6wlCNTs2sqJFfYtvuh9
tv7Kj4hQgs/88rhsIcpIHO3yX3btYxuq8DEo/fSdEZvkkM9zFQ+8/SOAER29fyOZ2r37BPYH3x+M
obyXZnloQJQ62gl76yxyAGPNFmnPjnHW+Z6zOLMESSdLoWZ7qyg+hECJv8kEUok1PPv6RXlFe4yJ
D77iAaJzVEXTLrT8On9DiNjDlJhrmPbloSEtShl3Onus88tVjy8vLr+bXU+CEA8t4Ohb+eMAJb7y
FGogQDrVmy/nqZtgn2jwW6E8p7+C6py9J1VDL2PzB9YRJoC2yDOqYgzTcAnnBn2aKL9upJmHxnQL
sS5CCoNmFReOTvOGh9v4XMcMQE5InpbWZHLJ1NYaJvtzMnaNz9NQXBYcY2saGkMdZg5KTC7L8WC3
jRyltRjl8egsLyg/00DwPrarQWm56NmWfUCDltpJfZY+zvW1EXHJ+HTOuTDmO+60f2GIhna0wsU7
lQSgOVPfMPdVB5GnETz/K+05iN60u71H6YvZRxorra6LOxDRiOlcsFbYwA5UW2Y6dDrS8Fv6FmLc
s6e34vzsNip8fIUP9JAoGU2fRkD7V0yXVRcrkzniCPcgTJ8sXHWbYihldQ+GKds6HKVB+DQiHb3g
D2+71QkydM1oAVf+9AELrOwrwJCR8ElGjm2bAWJ5cBWLX9FgAadP/IaJq8gpavuiZAoP1I0LFlKW
pYo23r7PDHVaWo2phpE0jgh130oaEJ/freMSJJnqHGYYkayw5AI8e2OQ3rlzkogCG03aowVesBLZ
uS3wriWvSrUvvSKCOV/A2jt3NRXEPuMzWl3BtWKNQh1fDwX7p2GntQW9mzy5G0pRLEd3s8WnRSEm
UdHsDura/YUf+HJQiQSggFy3hswb9ZAgo4FUdcCPubs+K86nC5842uaMfviRBCpX6ODoVhbW64Ry
6oZf8uh3+LDGV9eJ/6CDL1GB+BYmyGVGEqtPLVAVl74OOCfb4ivm73csAe+SXTsRqkuC9DoVF3VA
Zbo3aywJn7OD6qZBksYbFh9bnGu1Tzf/vTfROCWGO2ymqQfyJsUkDF9AtnqO98vnU44Mahr+L6zh
7gOJ7KD6WZfQAegnMT2xVqpAkOANM/Fj3uBu/qW95bBObuQa4GwzmWO8M8wWkcSUdrRh5H/IfEKh
bQfpfTH7bVNwKVI6b4Ju8B4Po2S/6t81gK71/QQ1gRovEQbsb6hiSGwvKDM65fQVs8miTIuhMbXQ
/VZG1AMpxDcfINnIjSluUGGX1Im8UKHE9hLR0+6HwEQP98XQ6xFs1Wmh7qj+HKu8E2lRTuGQ+tgs
Vl5A13nSlyUZpQWN2cqwfoJIhvoM5kaGKhlS2MmuVv9MJu/xtWJWTQu+dg54F4avj6JSCeV+/zdk
/vbHKoqxo7Dpp8d+DGqFz5hNONvBg3w/BYG89LeO+ZRem+8IEvgsfFRa5MQhzdeOkPJM20yV7Loq
0kSThTX2LVUNB8b3/lh4l+7CC5bh0eo4uauuJr70v/h8PsC7yFqtzysYnxWhdY/oahX6e8QZZt/1
aGS+Xte159fCWoPbwbwbOQZThD62qE2DnsMlP5HppLbToXnGCXOP0nGdm5quiL/kaYQcaCHiePF4
eRdkvWX/t7Cf0oSVRLUXp3X/+V5v4hh6oI+VFzuZboImcbZbOY5n3fPvfzueO9gOD6ht2IUIdmko
pS6k6FmapWjEB+3DNshtg6Wsl5/hAE6zOSlblyzsG0cznvL8R6Y0jrEiboPjodQVmpSkKutPp4k5
6AuWR3BjpJJR9vrYIvMe0Zf06TNfSbMgg6FOEtuc9vsHPK8YrfMrT8mZdX9CldS50yhFSa+76Hgv
bLHyMtkuBgCRvzb3zSNRz9IwECV0fy5qlC10nG36HYJmW/1VVWcsXSGuGnNI3BhXwpb4sfUYmZBU
TlBkouN/ibZPMKhXBL2c/WMFrxFukEJuoADOkJxy5HmFASNDnOKudZZXYv4OFwSm+bVhF1gevdtG
abHzWpq0wuY4QVsNPPKnTShtQXOCD3eWczpY6WUVVd+AEf/MA2GljRJ4BLRnJMQRK2mFJJ9AqglM
WsxPTEhu6yGGbDiBxTX6opoDR+ng+jjmH/Xe+R+hoQ5X2FX3YBBkexix6s/0rTKS/KMV/BMwGgAU
dKGYuhLHjZUp13qwRI4KmBCN4qhKgyo6jqjfeZFKDvLtB0YM0EEbkBLRYPia28iK41Bz5mJPUzJk
bwhUhvvqT/muEzK5G5syiW8sMAgoc/ZB5lGmKzJUwvyr/+rV6fBw7pGhxGUIX3fi8FkxqKDeWeOZ
20VTVR/Ifv/sHm+6uo7ROqxvOCdvowna3iyv4oON7vgIoHzLUMgRHl7pY0piKHXrNror4pa0S1B6
fki7Zvj/pfPZ+3bbLprh1bAtWP/bPv8J8TDwEv5VLqBlgpmNRSEjPJE2a0LyMoFhLGHMh7kcXubl
1oH7vpF/KsOj7VcW//2JGifHgDGvjzzjhTxu3zGDXuq+eFBTzCr8JrHUGs6BV1GuVGk4D1dG2Kza
m5cnyw9yC7iopD/D4qg8NOEMHLuOEQR9YehgzdM4bsbsOkkV08KbYvXz1LfmdjWuczwDn8G/G0GA
bH7mo7o9yDTio5TvE0aLJgRybLBnLKqTKZKL7XEdlLJ8F00HOIXQ/XscVdlEr7JV+CtCLmTu7NFb
vtKWifC5fQokk02pH0YMYDDJmIgFKINAkCJITaUV0I4nePbUjT87FVzKM67KjuBTR+kgBDTSBKsA
xpgN3c1hqjDyU4Hwearyki6SkvRXVYyenc0lBzCWUwxDz0qB+DFexhouLfHJQPayKZw7Pe2SNrnd
RZdtN92D2+Nzpnd5B+qEagHqd8AW0fGAPTa/wShI117Z/5liz8ThYui2x0Nq+0JpAKD91kInQv/s
XlywCKm6R7Z/GZks/vJhU198SvFEK9WFm8WrzI6I8efZyIedodhL8fH0Y/xPdMM0mn8VpvIkPr4u
C9kjyG9R0fZkn+8IxR2vzTfSsUWEKV6SKkfZcaPJsmTNo370O1+mewfdbx6oVliw44LnD0FTnBYc
11Jl4wTCw1QyVxr8c7Sa9Eylw4Gx/HNcKXrAG4N5Rzcumvq2U2XszzFtKe/bq0c5PgnyiBywWQXb
pjHvgSdVGh22bp1VjmP7pPLel5K6ckVG5qsL/nTz9bP9ZzVhlLwL3/OBl2WhegOSBWFiYMdu6yTv
bXCsS3+mddgoSXtPgz5fLyGRiZBU3Lbgp1WIgTMH85MmcR4/Lon3/NXHuFwMV/Vxm2tVA8FqXVLh
6HiN9ykx9OwbRCZfLN/73hke0PH85YzJFjAJCbN0MXAIJeADyKhN36tSRSZqBeQh4IU+cDpHq/QH
MQRLQBiApa+WoQvBjKs4Aclpk7SJE1gktN8B/v2jkRaclJGNc372LgZOQmtB2Xf5ff8D8iIv80r0
J0S1Dsy73AywHeQCnGgvWuRXw12VqisYUZFNrc953fVZHwgEuqXUoQ9aR+alfPTOziMIfYa3YxJC
EgzLzPv+zqztI2FrVeSCRj0bU8ZNwOjwvLWsX5CcaRkNKQLOzCU9Mjo9ZB90ZwK8x0vPbB83Tc4E
l/+VWCu922v2K2VbCrks56eUUPm20MQjLpu4xvRlqXI+OMLaoqKBzJd/W8+kvRVIeFbSh2LpsiBI
EwRfRBwCq74DnOmS29dENH3ENM/5eG2VQVX/v6JmOcD7O/Vt/vJ580eLzNFi4TxOhAPmjjF5kS2L
FiVxsKKotDYMt0d+/aPCTuAy+CYMogtQnfKnrqla/XVjIf7baZVhEenpvnIZLBu07APgI7aYWYgs
RyDnQ8dKTDDX7ZT6V6ErvzdooI5Ug8gSFZSJQbQWz8+GnE3TTaa1NrKOwL/Bqw6FVJ2e4O6sEwp4
aGydb+4+Fcvyy3KungQHC+Kivis4Q+dmkFY+ZFuI81tw3dMRKh2UOxsS1yLNJyvyeGhfeSouw0Kx
0A3bRqevWFEJ5WWcyDLpiegOqduC7fxTcPFNUgDlcwD58Q/WpereD5L02toH1XCRJJSMFLi9MOxZ
o079Z6mJKgSvODZnoRj9MXT12IhZu4KrSZDoOFCslGJHj5K8HvEBZyAzJ6i0ENhL8srUbWVWosI0
xFwFUBTjAL0X71K5ZdNEPrcfTZmZs1MHIdOOebAR5PwbaVAofncFAS4Sazk2+Hu6datsHTLx4aU7
uDFS10BqzyZK+O/As8uNoFhaFOphwv6bRxhzTTX0ks2J7h/WPFwsCtvQ/rp768kuMt1oCV7b0n/T
9WcJZSVBmaYdNYgdFMMaN6W+M03ikaOH/0X4zBkaEtP7C3p6p22PiolMjyHIWoAdxMvRhwNoV8LU
DQ/C7tNhBcFgDWbqBGxlyKvtTkBiE+mrbRAsvKJT5BsuJGn4IW5XIsVZD8E1yo3K62PbUSev1dri
dx/NDbBlCiUJtT539WBVGMVvYcHDJpvIwKlBd5M1svMwnVfAkeQqfyJdmH5gn7sIkJJhtuysgPNt
fyhgOnHoM9dqXqH8Tb7cUlSHeIKcrB8fSvY4+OdLBIg0TbJMFk+N1Jx0uu4J+gESZ4MUN2UJzUF3
O8pxGo6Z0G69513JuD2qpYQYHrnRrgZsIUft4CT06s2WFqGOmyjDUMHFoxWYubWbkMWsrPmpW+07
mq/4kupXrjujIFP3fN5Zejn62gKg9XdhWzQp3CEI+jw1LF2PKozhn25pXIaF81n7aUSNemKaJrRI
BY36GNJDh0eQnhfyvigquaddemxVLQcMlohdQS57pJmoXQlGvFCceQTLpLB7neGusT6J+kUxnJsC
1B8CN+exBmwnbUN5kRloDSjit999El94Y/93w+QLb9lRr6Xk1b0BDDpcD3AwxbSFhb7iwCCDBH2X
YprRMbYZW24t8aXbV2XOiJMXjbHQniYqrjOkKBEqgqoq3teazu61gEGgUtHFcV/Zekf83JGqDDaD
oUTql9/ccgjOyLiE1DC71srT4HARh+sL/bJ3KiR+Ld+WmTKfQ7Sv7r9WEPqL2dhLMaDlNY7ZOJSc
UJ+7IAmyUxfW88Y5IEPYzedCHhwbOwft4fG+kQDoSeMRIKz7Ofag66KQt9pcWMjQjmt+LaG9Jcgf
d30AdArt5jMDpjbG1PRkyVFk6WD4d0XnP0ZN39S2ceFCDKplBDOkaPag0rQPcoK9V9jQ/ihii92f
eILyaYtfURGbJWZ1QkDtNK/wjB3YNdM5g8dfDpqaTVgvgGACO/d+lWiRkYy2KvNHNrKN2FqQS9gn
eyyv5EQmuo58xwpyrAinCPRTw+9hiIYVi3ri4R62zjKipnRBT6us8koI173Bm3ymlI/mdqbfnWBP
5ruMS0G188C76nhSwREfUpR0cuqhmh6BiMySNDhYR+/PVFtqEa2Sk6mwRfv9QKIZJCHZUYU1HTKt
BBdfny/KVRMa8HXGcJ5H625YI5QNukXKPZ8vSD6GyxURJEllJIh4I1KqG8/7O3baTdSoyjQxkYn2
y4SOrMb2NQnWBQpqZVN2lWe8lnD0rj+AehiWIx01CwkGkP6k8p+Nkb2VG92DTK2JRG+ZaY5U6MiT
pOxVwor01bZZ/iKDoy1FNVK8KXH64CYLdHMmXLlupfQZMy3/3vNtxwjaRRVwTI1jHNscOq4+GHAi
8b80lC/eju+ONAkQ9hjw+y/mq81+KTuj8xfdIr0G2QShKM6rbOTwwPgM4FfCPl0TZ9nCGvkfm0Af
hnoTA9S08l7V0SmBSNB6cKbF6jZCBu0Onqdq+glpwelxLeAhSB+LSf7q/KdhwN4BGEQHmG/Onfs1
CfXCiRPtxmC9fYnVFLwa8LkyQL1YTH0eSTYtG2SXPpTjwKsKd+j2OPhlk7k/1tN4/f4pVXEFQGcU
tSQqGJsN8BT/2FKp5v3G4Tg8MSL0/LiqlcVvNg4Sthi13zs2iN5zGYOVC9tq9XyfGjH2brIhFYJI
CdB7YNFwXEADVS1CchWuRRzd6qozK4ky1uAZy4zEFBjJte1hO2VH6xQXzWoJdZXBCv8SiOMve00n
QTnfaFCqdkgP8wAZPftx3mWCZMkfakXL23xYqoV56NW1kHYShJjdz54tjO6yMB62zTONIVoGexLj
zzZUKzOs9Y75zLRbUAd1RkLICznmacEqPmHYOl5qcOYBliZHU3Cy1HAMCr9Ja4YsXF+2o5o9mhQt
7nAGeH/U5+LOAS4AtNj+56xWG/ENmrTT+ROiQjZM6OYImti0ZDdbvkCKOihQM8p6Fs74sIM5hWuu
8ooCDRNsJM0uVNEvy1hGYRfbW4wj2w9hNNdIaNOp23qaScPaBwDcyg6bzVKmXyyTZcFHc8qDmSV0
6A+Axyx4OBLPq1IpZfqbBk2axn+LGiCd4TZ+xNPWTvkokpisY66hotMf8iYplkO7MJKRx7FS8xla
ubAikmbv+HKkj6w6R96dxiNSujh7YxtxWYx1gZd5nQuHP7WzHjezkk2idp7m4RonUQXT7BkMaqw+
VnP6LxZ7ntEoFjyfJ/FVUkClxnwsGyMURRZPT7sLDKHOuMuPLMQSQxibeuMP3dd6FyeuS0TmKAkn
I3J7EbGc2Kymu1Xh2xXUUBi5JCTu1Ce86Vj7pD6wH9qq0Ls8CFeL6Cd4779gjTeYAU36Xjt1F0Xm
rOpKve6f/Nl1KhJa5/cmWowDxE3j+yf2YwHPhIbAMxvCeVQ9pFrcdSqyHvIaliEJHHQXLEEBILZY
g+3Zx4e1Q1m7KiMXHJ7UjJHL6MHwUPmLG1fJmvfTs8WA9V+4odl+Y1hc+vznvU7qnXRqx0yE597b
Mr2UjU7azEoWCBCAv4P0/WeUaM++4GfHHYbh2MG2w6D/FEWY5ATsppOO294mtDF+OqJlgh+UPlXQ
tmKWORenQ6bA1OgvYfrx4ZbRAA/FEI6q1Ioly4/40UayaimHq5hm1AOTU1PKjqxpb6T9/9qTbvDI
ybzicHHib9CW2U+xPHwes8kzrT8wjrhAeZTLEJFLTnueVG/b2pHIMvtu40gfIZTqtwVuojZeHQXX
yxikJlqDjcnz2aSIzqygid5KtCoC9zGih4OlfvuPvmnVF7Qbn9VxsynMS12pBbNnx4/wFDAEuLNm
8HLuKFqqXoL+mEvFt64EfxL9aTn8R3jC4MUJJ+JiQ6gvLqMrXe0HvSJ/eBIRQdghBNPC/GS/vOYR
bSFKvsYVRpnP6zMhb5AfEXp4ZZ9DIQi7cMyR1fILt/94rdhvOJeDsV6qoE25EySjGyd4IxvgBy6x
vurgAdoQSRDn2uTsE2NtuLo72D/M6ZWmEpqn5rmFhbaui32tmnZPl896ExKioEkcNkyPWgwCa+FZ
N5AYwDAwZBJ8rpatHiulnnFg4KfHp+e+h7Cu2YLzcXvdU6LoXmzWm2rMt1FcYpONPRpuv2dhAP5r
8Ck7Zkj37aZOt1hbnfHHTfEJjpu8CN3IDHW83IHOBE2MFoiXvr97oF7m24jpeBs9y47nOnbrYqq/
dkPJJOwu1cIJvR1ntvhFzXg46EPgrd5BPszWx4nY6Takx4wfYT2ONHz+giAAF5SOJFFCKT6WnAgk
4Ts18JY9E2Pb1zWwBomM3ifD97nXN+LcRfCUB/AQ8ZL1RbO31wS7xsPEcVMqePMknbrXUWz5ZXPE
7OmJy9/c4mphMnAGUEDKpWGxuRVPbip0vSbNgX7GJlkdZ/4/Mf37QgnYs9FatNMN8y9m8QN60F8z
8orsA7Y6kX0f7Ymxrk7FC20p0PYH/mJgxccBqQ3+fiLM6fdo2e7aN2NkOo0cq2ql/81sHDcJRYc9
1kHc3L0HGlvucndnsI4UEkN1HR4SK0Qb2vfxkREdk1htnbs07x9tA7oUkYf11srdOCnzVJ5BzLQ1
vuC2jQ9cUqpNHg5G8xEnXpzvKweMMGbKIHxYFPsl4URQj3jMY11KqAs9c9349ABKiBzaQlZtiKhG
lKQ+IVqQLqBU/j8awKGGqBYVtz84UXxYBwZwYehsWc3Hk1YIADmQcy3CrLIO86rscf4YtDePGnZK
t3wNmYlXmSyYhldHuoL+5Dxuh0aoliFi9d1QrViPdBl5hcN44D8TnfwG+BWIDy5fBxLeuR3artc/
LyhZz6/TOlNnQYgQFJxEEDERGrAysztV6YNqDy+Md2pEBodnA5D1dTRZjCb0EcU8vOBLGiZHzGq5
D03AQw4VcNnAiX3tDe/NyrSqt/w2wiMQHJjgAXExjYQ7H9YpbxFSXhVqwB2kVeBozAis59WM5YKM
jEm7j8TevIWgUE09H+wCSIet8aVPpfuNSxUy0VSoLsr65YuwPfz5M6T2rWiXLlulAY83mrbE3mhD
vJrg9PjuozHwPktLeChxNl80JU+5quNtAPBPc4pbH61N4u7n2pAeiO0fnmdtXQY8cKfJCMIRIXL1
MyqN7EpTr6sivHeBcO/kRaMCNvWvT0gsDcgHeyP+4tprf8jSEYzrOeuhnwM4GAQONQHswBTYI9dg
LS+yEkNnfvbebMYJFmfezHWGNMqBgEOYvelAMfzuIS0CXHybN03ONoUAHXJ2R+R+Twihy6rtW3uu
sXELh3DLtlRnDzLabQVwOs288THrYcSx7kmwa6Yxu9FnYUZXpeagAAuLPFxY0F1gnim3IUOPyyvC
muLWoRAYg6RRWAsJCNSbutKLnDd4DJXCvcgAGM3Bw6GA4rrMbKJ1lmpptyZtUIoNWfNNg1dlYD+v
rTl0IK4AQTTME28/sJtOFYkRt3yF2NpHIs2mpwZPg1wkBhWS48rdiNBO8/teqSg6kqFFzIHT2dNN
PXaZT0ojCcKaZI4w1aMIdiqhLmMXU9kibFygXVkTCmZcWtiIQwTP57X4bUbUr9j4digbyt/QuSq8
yUUk4qOj4TmO7DKasHosoFRDne1WV4ZcpDupcnWQFB/hIWoNxRyqE+2NmSYFI7Lfw5Cc8H7S0/1r
aRinaH0h7CLeZCMUnhpKy21PrYgOFQ7GrFlkDUtI/ZDUuhXBDkl6nGmjvEUQMN24k5F6VF/+lVPi
Xi0unlrDF345lwIpCNHXex5ZgEvBsdzyzIMhek09Y7qpYUmSmzwaMqJvjIdGiJ0TDgbihplHLTAd
m1IBIrBwQBSQwajHzRpG31Imjq4ZgHW9tLFNkVZ94EeMtLvI2AgbcHpjVQDgNw661P/7TDbKUdEb
GBSPZ7u8iCv0PPXo+0p1QlhaKkqOzLOkFQoPAiu2LG4sf7kwanOh8P5DwKy3NGP65UATKsCcE9Bg
Qpto5KLP0xkIX0z2p2Q3v2Ek6JBHHVkNaaHvCGnKiPLvXF2+ppc29i3wtjGrow+QYceLn20LqkL3
9+KghDDZs609Ja/QnDhQCLlXWGlzVV1BJqFIDr0v7LSV+AmC1DlZqnrjEZZLXpGwg7ujzXrHZdtL
sLGKSlIpkUVg0mpSDuJ95CxejLlKlEDeIEMGWaVq16s9B4/sGJpaIl4HbXXXSkVs8OYE1qeg5TRu
wupHRhJ/rQwJ/P8q1GFNmDdUzpbGXmjCX6ovtipw0LCO8Mdj5LpQB7bmeNlHY11L4I7eQJJFBlic
yrfzIsi891vRL3/8Pu48MJn2odPF0uIlBTOfV/YnfydxpMopo5VSCxkNQndF/ECOAvdvwkxU0iPn
ZPJLUY+7xM5jP4MLf2+3ukgIzePhabYsN6Lyu8R4UrDitin1cjY1s5TZuc8M8vEmfQbh9qTfHbG2
WKmApNGGdSjywTng4DF2wXOL1y2h8nJpulUdcpXA/2DPtE83cIzzFyHiwNN3SgaCDiUHKelwljHH
6WZIGUeFE2SOKiI2FdW8+0OW7OXh5+6sY5T4c6+8pDrtOJf/TFzohr18fa/0bjwQ4NEpMm5UzF/C
S1f31UgnQSo4bgOYUeRVwmwn+E3JXHg1dZnrC1Mj/W4lOwF2lNRqf2vBk62uuuZ/LVUWQmlBfbw1
IoJvHAp/AJWAktG+NKR/6ZBQYtvBuYvDgEZzvaxxI7VaKd+P/y+e1Q7hrlNm4Bb0AKomoaLLERry
LGNfOD2RoPujs/toj85lIDeGAoOa3IZEAnuqDBiv99AY5K5C90raNgHJ+apE1lOiY8NVYSVD7C5L
yR2tt6H9Q/V7r+TBUV5YEJTJ0xhBIVKyQfV3t1mdLLZtqnUrOgYmFeD4RJSnIt4v2M/wq7SRUKjD
hdNfhujoe5pXIMtxOfopZ4OYrEQ+1uqIXO6vFvUv3Z076ePeBU7HRqkadBH/I12e6GFrdRAkRb4D
8R3Jz+SR+hvyjbGeZSziXSjhWBP2JColflZYwrDkYoropq6nHYqqxgHrjxgV7YVymckqEHoqrmdF
g3yZkSr4TDCfcoO/NahmGGJe1T3/x01LNTNFdJS+nlnG1rbYNdocY4kImJqwjjolzOZccy4FKVM9
tHlLCbGYLN/jE2bKtI44qgqToboQDHB5oCxCuuGFCPIWCnZrFt5GNagXRXMQftwMKiXEPNJdOziJ
tSeoSXbzYVfyTRA9pc40NtT3yK/OSwE2YtsaKZo7IPENKZL3Kva5i54NHIvEMrfvJz9ZZ3pOR+1r
IK3wkO7H7FiRJdmNUJCZKcWQV0to+DlTrvywJ+vx2CGKNE2Tri1BBfjLcFDSwhYnuGP+6QpEz9LD
2esl5hxovxbVhGgDV/pZu+H4rowVtnvlbwq10WPBZBKn6U0owHW+JwGx6WH1ppIdh3Zw1OLOVKE1
zAhvD5GMhw9/e+MdA8mK+Dl0TQr6Jzrv2kRT/jNFaI8v4Ve1PnEN/poMIzFumFYJxJh3kp2DMm6M
yc/zY17GlQ+aMMiLEeTMG6T/sbTTLMqK2JwYWxclnOCHSFFEW/vQ68Et9/d8mqGlMLOMA2xVAwxR
lfzn72Sjist4xBclZ43FB+/Asn4sMiTvfNryCOsRnD83N7CdDPgfFuNJojh6AwFcvIoF1EKlkmDX
Yi+V2u02/LFnPJlUXyEtZqsMnOtVEtNyvzzSEIn+G82Vrt55Wxn/EAh3sesgkWF9jqct3AOf0FYN
KCY8+qq5qqtV61WAEyk+HAyzzUCVGx9F/3xvlgCvoZOjGayEvabs3BC6e8vaVt1uzHl/V/7tEMlO
uUfKLmH9JGmSpusV4XeIAw3tZmwWf7bhIVdlklu2Ackg16pVTiUH3zgrqym9A1clPMA3qkdJb617
CQZoxS9Lph73oth20GzuJOrShHADq02EQTMLAWEY3kkxGMSS12KJ8JkyPCRT+yk2yNsTGKkfaERf
YxAIJh2VOw3Zjz9SbxM+MOs85fDS4/tTyXKd2874v0ptO4GsQ+79BKZ6hnb6+NH1LFdVgL2o8LpM
VncOy40+Pu1reD434M4XC4nJVa0/J9C7a8BT+GOmO5j59FJl9kFFPt5ejfU4BQqw3s2K1KOiMHmE
xzHx8OvMoPvvUjLLdFdM6If1XxaBd9l623NP/WxLkpDFWqLPgitvR0gtuIsXePNKK2JnOUH5jc0/
CUy0JZXnrBZuOFlgWWU6Zm9O8BRrJTp6cPkninxdD24teEsxsRU4uimhCAJHNR/xWkrTDnq2Kd9/
gQ29tVqwYQHxempFLhOgWAtSsf636GdU0x0xRc5h41MhzFrmEvunWRW1eBM8w48DMhTThvQHv35e
8Ijrc8rhJWCxikZzWGbNLX8c60IXbOD9NoZ0+rUrX8pAp3m7i4Fx8gn1wuArcBEd+ZK/Vygjwf0h
MFWgcfnDZ+V2G2nJ8Fjet69keXMZHRQFVsM28nzaoWpff0d3sS9fZpDQiGJckSHrv2EU/iZHICqU
pVI0Xl3fnUwwgsrTWzZQVa6BwiI6C/IgfRKHpBp+ezK2Cp9FajPeVuL8DSnYZxt3yF/eG0PTUODi
7r0PAN69Fh4rCdRuHTU4GgziYF3dBEhLSADzJHE5DB26dEXo1SF3AacfcY/u7n9IYSehmW3I3FIQ
i7OwFDcGHDxb/Zz+xCHiC9Vh/NRULdsBOKwoehD4/BBLxRHUpwKn7zjsOoKBxoN12kz7Oemuxn1y
GX5b1EgJVtaR/KA/Qb+msRw0OIvkawXPzuwlHQEv44weiWgqsBgVPrMNiTqOuGBCtPhyCAtXwXyY
d/7FOkJQh+R6QlwOXegEXzRD5C3e/cUDJEZYo135H/yextCXXG4eyDFeKhk4kpCa3nZBxstJRQnv
TwfqEze4+YkIGyo3g34H86fX6XwlG6slVvYXFTv/o7GKS3EdCGaWu3+iFcozobbX2hlxbuY4V5eA
PHxWCbShzTKyZshAQ2JS65oFY4ChoBzB255zp9Yqa++04kKIkVsWYAt5oB7cU2cK26GIIKlNd+Qm
4H0Qg4BZS79dp7Jl5YwkZY5OYq1slzbdqmFPQsuoxXxL+fkvswZKYiFrHNBPtMjLyjPTNvwn6s35
Yp8QK7tWqoHOWQ6UOYxaD7unidZJamho5TAoeCFokmlMGrodlgPEeqL7jNyHdqQQ5BXUBFEZlKl/
GV2YsoGPXVnJgfVhFuoGiSGEG39nMXCRrnjb0X1Tc7sUPH/wX6xAw8DrXYjBAeCWUHAe27BCxJ1X
L3iKbHvKo5RHprR6Jk+qkjSV2Y+zgeDN+KyNGYr8w6vdWgCFMnPorCozl3nYZTK/92ae30fZJkkt
o6Idj4woSqr2vD4mnxfbTp6w4dK7SHc1dOLiL5bxBQL/QCM5uknM9QgTHqLL/alEgp+Ktus8jn24
gglBNazueHyC9I0sg8FZXuR6YJ+Ag+zSAhM3dAQkj2BKoK61OsDOb3Z6/kuIukc/oP3HL0yP+CVv
96vaR+rvJ3BUggZEU/1ZfZsvnVcJ02VnkivMIkuFNRqHFJXkhHv/4d9+gW5cb9vn6ryhzRDkU/df
gCKd+zMdyo17lF54i0gGrBw8CY056Oh2RlK1LJN7RkNvcni3+ldEI/OHHtE093sglw6ibrDhZcQd
dMn9d5G35JaVdEKsN0MUHY7Y58Rs7/MIsY7WYNeJJJxV0G03x0DzBDqX/pmWu7y/znupMT+Q5cH9
A9KOZORVwVPxqGTymlCFpD81eGmHIz1qeTs8IE0LZNEDBMtrA9od8VWG14R7oBfCdhRD2/gk+B19
pYL4OYYosiOOfsMJ4Uiqpf05+3S72ynQ+uA6FITVLbXH1OYDCflxpQA6wswKccwVpOjXSeZFm8pW
HYwTLMxmhXgvnGBTsq1pf+Yqk1T/gggCZ0D8j3IYJ5izKHOBAPwJXq1YC4kVzv9twXZCgkCgYWGd
/2PLtLnhAsaYGmII6ln6krNUc9tztuordhHgmyNdMkGY07F0QXj0KvOJ1nGPj0CHZVKEMWlHBCIR
Ki5NR/SdmPgdOEYnuvzKk1Jj6QkZnbr5sqvEaZ0I3iuZFz8e4kvcpx/+TSRncrriQ0QtnnsoGzDJ
qBcY/SQY8LFk+XF9+we1CNTfKUbRgOfwNZz1EzCehIqz9psb86uS7JFZIwt3RgxehaeS65ytQPvN
iMWc5Ilt3CCbEkSMEIXLWm3HDrQk+c3wkG0TiNKxtIGm4JCe907TryKehlx5UExvm1HXqFqhP33g
d2TB56lUvR3s85VQF67TMxNJw3M9tpdo666m35lsAMdO+BbJyIUsh7yFY1Kl946QByexRmobe+Tg
ci+JsraQYoX3/e4cVqAG7MNIOvdJOKF/WzgebAj3m/UfC79+6FMARzGCAL8WT67AO9otPFdSoYCA
qV1fmz7R3zeojZIIuHAZnxnuLNoD1vqnZeIVgqmgx26XcbJpP1Paar1z6z+y3lNW+ibArtlqIWFS
iD7JfxteSSzX/cZz9KRa+VjpDG171FYoxbzaswSewhznmGFfHmi98fnP6HmYRGFevfpkFijDSCFx
Hpj5+iDsVdEMlal46z97aU6GoPqPRuHEOy2KHqsA06/4/BRjf7bFZrUA8NeU1OuODWfSnaeqSlL5
2umL4BxS7rizbiBnj6cVXfU31EPEaH79NAfy0ZjR3m/EBq7eWe31Jb1CDXyd2CqEsHbWz4EM87Yv
DFYM9/FG1iZZpmA800aGbXVs+7T8QFUPsbKIMvKLbn8sKsFcUo9W3Wk4Q4aN7cMfpgN/nXdGneKe
r60JixuNR/F1o3/JE9S0C630j5hBs1JVbe/2qhkEd9rKFyvGmWVSPwjNkXQTxJJMYPoE6je2cCQx
ym66is6w+tMNB4jroEc2qx6C79TEoRHwciC/cFZQnlWVukHqyqOt/EdUK3VkIrkfQEFuYbCtDPcc
dmVHytUhLT29bLL4WQPrfFbZg5oSdl3JDhMKJJXmxuBxx6jOJvWEUNHpOy3j3Rm4fQdvOLixpzuq
wb8rYrJOtOhoCspblEGYwjjP821rusBlYpNvBMqcz6MwuJwQ4DX+hP/KPZsTDma6ZSJJiSy+sy09
I+Vh8gwWtqLoQR2wUEvp36G55WlSOa0jIsGVVrGgPctvOpaPN/DTRGUKwndhPt607fwWXEb49GFs
m/tFIcSbJcF9MRV3Fx86PwIta7kpDjoVSh1ZEGg1xCAZPcQn6EOCxci/PVhbIr1Kp9VLgDt3xHD1
dpkSCmSPE9bgghzwpADwpwhmtucmKWJQt4ss31YM7Fi+FKTBmwaxj/vi5exvs7HeKgxhWZZfVU57
J0IDhuOH4biQd/NUm8pzMIQOgJtktrQP6iZ/4+fd5Kn5/uupTWNpR5cf58zr6nXmTZN8F+nUJwhm
2dfgN9kjIqcqsduAD1tygTrfL7mtqNUMMUov/8WDv6l4xsBkzVS/Q24dClPefFA7UVtPdUjLrCuE
CD+W2yuGEDIDByrsosoV1Of2eTWHAP5UvGu1atVgDNPxAUyaAvI+vGm5kdWOMCRXnKQ8Od6eeAia
otpMb/JXYXwaGQbEKcyJDFdTt4k1vStQG1RDkICg/g2yOUgPSjD9zRIKYqIfHH1InZnhQuXTu9y5
w8vU5R2GPFnm4s82+XLuAdfaUowB6zC0uxlu3v4eEpuYSEsjkhK4Sv9MM8J4OgqBWC6d7oUsF4AV
ko3nWPN0U+W4cAZNie8iihzhyWrd035lKypN/3cNPr8M7tc302BFKK8u4TEUaJa+dYl4S4npjkoW
DiAzsUuwIxUF417QSiegwVuj0f3J+wQQeYyxQOJ0TojdlUetaOnirid0gHzVN6erg322tYm9qwrf
ZNpPwc0uYPpFwpZVwiOxiQswBTn4DMDzSZdioVyAvDrkRrTYQuBKBYrmYZ5VC4txRJRTNrk86O3d
5ykNSSCvdHxK8UL1dXX+NzS7S1wGAZ2rI8Z/fc41fBsVlz8SNbXbk1VbiyVEDtfafYknxTUdWEMy
7vH/LURGiQ050sZc3rbm004skLprMRHYDXNk1Zn6FvEOVMc4VqU/VPCii3aiWucZd+ZXB+DplfVk
2UZXPEcqAPFTB0pNiKwxmHyvBD1eoJmoHm5xvsLUK7rsgAH/My2sSszo8SjYeRl4pr2OHASrBWo6
t1PHZbP3NPrlMnssmVPPDZpEyWpZIETjNd5c4Kz9dUI6F8G5h/4wsKcS2AJ5nV6qZvOJua1K/BSL
qu2ufbB8YOTzKB30Cmw+i0jBa0GJKD54cIF13e5r4QGiTQ5WqPPENib7ltAu6n4dElcZ1CzULj1P
DTHi23Uf7SF+/3X2mYXIoz++INilj2nyKcJo1wY5K2XhDz+WXZQIs8S3JlaOCqKp6sfDaP4pp+9m
0pVH1dYx8Iu5pH7LUiFpkK6bsRDvQhMBj0bEhUkmnUA6E7m4Qo96TPzavrQ7J/qYPOzqPAsL7iYf
tXyMEPv8xhMY189X/iERFDsm1Z37SZQ/6eYb34USQfRH+FhLUcvbQF0f0GNzn2LyKSwgCDMYhri+
4dWwwOXevWExMAVKcUNX18vL74PHBYFVZAiMwMr67bpM37ZtqUePLGw4/c9+TvPlBq5we7eF+nHp
7ZqBmoYdR/4ALLsbXLZFSJbEUskm71U1/jkZKlHEH4ePBui6+/Ybc4wq+LrT4QyRVFqfWtjFbzLa
gSDbUKi1nXYaYOUvEhcv9ZEuRrXJhaWmb1PWlJvAWtIRgwIQxwhSiDUKsT7zhKpRBpMV6LLmOJX0
dJoH3Zrf3P47EKovEY+1aCNnpJdD/3QY39vw+Jkh2HBYiu5h5UUa8XkZYdBSfza2pGSzo7ZY+qgx
h6u7zfptdUS9f0HJEAXOHaPyrInHB84ZOZDmFXQsT8yGfwFasadWBbGDnOJMcH9jq8GtCoDDCBnB
Xy0GF1qOUybeC/PJ12tI2XoJDxxrdiJeCZ0gOEHcFJ8++RuuJ7CHyzi7FnENtM23OQhewMQIAjQL
sQZb2y70HvIum5RFMyX/G5YHXtJDIkvLMiPmpTAWp4iBCc27Hq7EW84DMseIu6TcnxkuJ6m+RGg3
w7+zNeLX4PgqhUxd+7FAFTzBb5rfcQKNXzH7G/DDsrPvNxGEvJHq6F+0sTK3229J+LtOB0Hhd+z4
Mi1rL+8BbhEnKH/Ub2KUxaLDZ3AE5yhU1oRTo9S7p5tJkG6d7XdRSywI5l9FEgEiOxN/Xwm8KhNd
DN2NI6pCkQ7VKpKAKCMy9UL2ho86vRt0IRw27MiyZzSaP0YaPp5TwsFrwTtLnBfP8z9TFuTTf5H6
HmUhaxJc4b6fCnblya2YjfyY4KyiajQMczPy7AavthOoo2IVOq25xd94D5AtXkYAPfadpg0qhTw8
YGBmWCkRXaTu+gu4D06mdadbI1K3FHRbJxIOHLl3y0wrqNZWuVfoSluGPMANpJRRQS0eH87rz42K
No1R4s1IPzb/DNL3aX1gycmjXeB0UBtI0h7+ov+gRs6UIbNP3a1dlReQb0gBw+U66OigGSQse3cc
7Fgo+V9g5OMpaWYWaQRSD02nATOQqwmPDdPWAmJlCjYQk+01WGhnJRIxHQIRHg5pz5V5ckq7y2Ze
sl0Hg/9ntnw2FylWPMneV8hydp2Iqjygmj68D45h3UMvOxxKRkLvORIy8/V/p1ViBwcwtJ2NjoNx
ldyzWFiqMKOadeDljT0DeS+BjIjAPqBCsqU9Lng9g4xJcFz5v784YKxBxabRI72lkIKUD06XC3AM
gpY4H7RrkSUpO8NW4uc+uAMOJg3D3XLLAlQWB1R5t7EF61ED8A0N0sX+ERhtg0OZUoQL0NYFHPhn
71R1StLdsVqs7jrFB59nrrdmoexVwLn35A7TMXIHAxLtM3KKb76f4T8vjU7xqe4bO6R4FXz8ApOU
W0gmE5dx7+K2VeE26QmHpw9QUSpyPzVLFH3WED3p4OBQFJrQ2ovqJk5e7JwXcyA/Q75aFk1xKC2f
VBUr0gVwyzKnf+3n5SJiM9+GU87/e5TAsZpBzqiXOMIjE/UwxKFPFs0yIwqN8T0fCWOxxTvc1pVX
wmvBpZr8COgl1witzLIm8jmc7oTY6R+LjprdNMDuHGtT/z2jP+DUj8KgEPbAgeHp7/qzeQlNDYOT
fQi+KZ9bGJXuYk3iBye9o2AFTl+EuZvm3bu5mqes5w7fxD+EN0LaG89YaGdUdVxfcuyxxFBqmoS9
6NrtK293JfCl094sK5/ZvIwlCHjWXE2iQYvnKetXg/5+YA4CVLB/4PkSrYnAHpmNMCaHOUBwCQF5
WKJQ3arZcTWVGtueB5srVYkZFpotkJK0Tzs2ynbTMx5lh02Dqxy6TqI6n0hoVJpDdNDbreil2kxP
V8pnD5nVGy0Jxfff/frGA5LaXH+b79R7jwcpeKOLMZ/15rAq8Igm+cYp7Qi7PX9GCJlaAS7pz+IZ
2fW/WeH3AjMkzEVML4U0DqKqzWKGZDfYMCm+O8ECjTlNSGBCCvoNX182WGSQeneaRfmKBhCiN7Km
mJsXATOx0BfDzoIwVAn++RrhvPLSZMFVL41SWVl3NVue+Zcgn1rW2ERmudN8o2TIMbjflj+Ez7MX
N0uxDYYI06B78Rfa9cLxw+lcqAiKYzDTFwz4+rL7Lggw+NpSj1iLxT5gBqCdG9enigXxD2/KhYJ9
2Cv89ASo7i9zrZs0x7dVMLLCl+cLGdr3FXPAi9Y6WNeLqMFiAWssBWQfVn+VFIuGRpf9duZdshH2
M3YHZoyWviR/OzZ1LKPx+iiqOwKVYUbNm3F2m7YxbNOjx0FPRsU/7zbnl+kgya0l/lHKyaMehHaD
Vr0OpFg6JP17klWd5KMZAfdD8S5ONA42EJoGDaNdscEN7bHCZzN5ZQO6nMy033mDC4yUS2WpIuH3
GfeaxkUsEDgQM4FIesl0lP86B6eW3nffoBgaIT2bII0bOT6TFI8OVRmiQgNfgEG+26o5V0Sr6m0z
Gc6BqDBG/GKiKdJ+4ujYJwiVlIX5mq7jgBWUwuWF6BO8HzXO6wD4KaUP1N3OtiLCAER51S/RNJbL
dueWcvASQwePUGQg/IaRRQTarxUYNpoHPCMMSXYlyGu5q9+8Ne/O/qOXBhJEidGBErjX9cwVj8z8
Y7s3yemmDPl/sfqSgyLH9hyzPUOxkJ/en1Qlc0nLSrvhCQWtBDAtb0oP9lggSwYyNvAmlcv/UP9g
el63RyFp+iZKIjbjz3rin2tYZxzYK9+jvwJFN2SsdbbReg5IzeECCJ+Hk5bzXAq5lf37os8+Rddh
Qq5hxsQVfP9j33+s1lSf0vpsa9vDApthH5z1bpGT/j0wDaQ3A6I4SPT6JACPx16b50jWeWMLNHzS
Ei1L2wJh+dtYeF+KKLBW7cgyeTgK9NrW7bhJ9mVXh5P+EcxIcYGr+HrFPU6oEkO3C49DT6XLulXx
cZcJBrDbo3LuFEBH43QHikqIR0LQcs0Ydd1p4ypsxL+cokAmKjt9B45PoP9mFzyvvNTy/CoitQbq
DSxFNcwelB/7ybcsosdVqJl5V8ncQ8ez0hXFZRHhzU6X+IQ6DYKUC8YnAi/VE4ODFwfAsSaykdx+
RN3Lyv//soaYCShP40Tri7LKtV1Kzd032sSRc3lLhc+XbvshJouBf/m/wbSebR5hNCRGI5isOJse
tnxTyfUzpUf6Oea2XnmZY2v2MHzYvSWJ4CgQ4OYzNVl12J7Busqq338X2dLgY1Rl+Fu7+srCAEli
L+PshzKQDoCwxybx/e1b0V5N9aLin3bZl9mNJ9tTJRfhBmiAH3LjeV5hxm0OoKsTexRWo5M1NX7Y
dvo19vIl3hl9f/AbM5xsMCo0WkxK6KGxKiBQk+ldYfVe+H4X9q2uza97Lbe3MRr3AgmmKJ5Ov0h2
GMJ2u9C0p+RAG2BPAYXSZZLwCV3DT7OOuNSkUPpJXfG54/tXGtIKRjnsxpjAKNpcp8j9Bzv8BZtH
aqVK35GgjhaUXWYRF06SwAMnNaTV6HhqXw1ZhPfUcIno85eojtG2QriMOdjhMtWS7PrP+U9xSLWz
R1qIQEwpsUti/PYr0jJpbDSry83bqHU5WKQoZR9AuDHFMr27r3nQc7PYJW2acpY84hnl/vtf9LY3
mEmWZogDeDANjEgs1yH9zl7wl44P5KKq1jq3yhR5nhZOWIdUK8TR0TvneqjZ9GOaK6aJG9VZ26pX
QM78Rbf95/zRbm4dKYBAnVagAmU2zPWhOoVPPM/S4bxDVjEBBcGhKtGIej9ZMZXW+hQoGWu76L0R
QpW3cjsciyr9HGFr875/QPVw/HuUzxnXDo5b/xiI6pg7i5xzstt4eiXh4uZcsQ/DmRT5uBQ2ljR5
ldY8dKVI4G+qqM6JGul801nr23qdLf3kRkUtdHcdERCNpmqohB3V8xwbm1UWWRHFAkOwUJBFHcZg
gwLS+LxLaMZCZvlKLQM2jC6tuBCC5LrXK6yHwtD4naPa3K2UXWxMxQVgZTe0HTLmAIR97mI/qqsv
A4MzCX7cNfyNijLxshxV1WMImNL9UZMrfxpUras52i+SdAcVsgLOENHvruviyfbB9J5ge669iltL
mKQL6QBo1QqC9+1BvFS2Onu7sMJ4Megs9jgTR3JpgMnhhw7OvrTBIPu4ccEmoam9P5tUWKkhwgJi
52wqMw+Gcc2QndpkQjEFLG5XpXpWVLBSNq9UjuY8ojE5D5t4gis+GLU84n9A4lOTOjvp5q81Uly7
n3OQnJjO5+orXNcKXz0tTdKrnWN8PF4SyPn9vCNaZ5g6wq/rz3xyATV59nIxuHu7vfaBsdVQcOCq
KuaXbwWGGVpmxZj2KITjOjJhcJgvWPxBAm0vf+LRcayc9RQfLc1ecFcpUwKsTP0N4FBuGmHeeChN
WO/J/iyxbV8UtA9E8vhlh1ESe0cCiOAQsbDr1G40JxE/5ouGN3NqAwYIQvKyRtp2dwBfEh0JW88/
YV+5R6cSgnOdkOiJYoJm/jDQ4KFqWQUWsm2iHwhNzjyUPVV7tKzK/BL2lq9/hsTonBCs/Iq1QpVX
4IjNkgLqZfNvY8IujYhJrp22bVsM8wgBgu8Dl+GNqtb/5XloC25yROupr/ZigVJfxuyAzMdFgba0
Is6A/b3VodX59JQSE97+iopAMN3FVVbv/LhbtM1yFvJ0iz5eVkYlCAotFBMtQ9TvPUeP84QybTZO
AecjfTVJ0f8Pf/fWghOY1lmdeWY0Qpi28//LqR2IM3DgQCj7Lfki/MGJNdxeo4MLx3qBgS4zvcnr
T9XPVBnKerAXKJ1oPdcu6OpwhgW60CzEiUVqdlXvO5CxiS7sPHzmkif5EA7JmcM5NmYszAtoxtP3
okpt4EEI0k8S1A4GMvzQe0Ga9PLXtU3aBmCoRmmjHl4Ol0IgTPG/2ryaHlhG9MPYJp84964K1nrC
62e6FLK/kT2+T8LxE5tCu6GeNH9TLHTtK6gmu/T07RktLeMVB85CieXW+a/tTdSKksOSDWu97wVZ
kmjeOqQbwFUL6ChkEEtE/CQzuBohpGVhTS4aKSxulg1QzEdB+WpZjPYsMHdCKt8RDarlJ+jJh8+7
3jf8G3o91JeXEvol4DZiwrErALNgfXZQlI1Hc4Mt+uHXBNsgjH380PyNny/m9lR50v/u5no/gZwf
zJ5zN+EKSl/TBFXU+WbuKW1vMb6+rqfE1XM2X7J/uo64Y41Tyw1E8d0Fm8pWfAiPe7+emxsWT+n8
Ggh3xtLp5ymZ5WJos+nciXwABeWtK7V1Qm5oOe+drxNM5+TA8iRFUQgnVUsEbQHuEmiwXVo35OwT
OYPOJVk5Yn4M9t6nPxEuNzs+/I/zHICDhPUo0k2w+RMwEKP0dNBUqEXwsVkmvOxE33zNkGbOoPek
FE2uuZMugsGnZohScfwfeKH58/eABT2fg9XZjF4Hi+oJAYb0wxk3497Y1imHwg6gzNNyDo7t33Sn
v/5R8IkqOmoa8zSHGuXRHx/hPdlfdM2Sn/tjfLixsEMfFL1cuRBYeguZOIyWAbFCla3j77I4uxJp
ugKedixuNRD9blVlqedJzVJle5LyCwB4y1YjubMnYlHgcpcdW+YX3p+c6KOknpgGT3BE1UnCuj9P
oRI/MTP5ewyun6mJirlol17o6BKJbIBDaEsVsUXFdpG+nsukGIXcPfok4DHYEH9f8P65LmlaGMTF
c96DQEb+sz957tC0OPaRV0u7fmqoDGAdscYlPyPAi/tjobfWtAyvkGrq73dyG0APpwkd6AapcX5A
wLhdY7RExfPmltwU8V3qMHp4TEVbNuKG5g59CpBbaV+rycajuf8bOduqKWQb09Ny+ddjgMdH7xa5
t2N6UOKtTKaLbcFXgDQ9kP4VBlOdUoCaSDBGZepIfETxDeb6x3RtMKwJBAx9a/HU+phH+kDzpPG2
J1zRJJ66JrEitN9Xg0Txp0RWlQYEXPWk3knRB9cZGbBp99JMcHx6nanOJBtC6rJpkuBvTOfDO1Me
6m/WL4pPzsMeHDNB+ZQzKcRU6CsdXNRLVdnltQd74MMWcgWEB9FfEZZpArvTIRnxqtwHN+YQOBhd
I0IrTGH9x7448SskIgDvsnjiL6ARmuC3ogmXYfcQ0X3N/EFe9Zlnc/Pc6BypTrs9fA119gLFXV1x
EBOsh0zNeOAWuvB2nV4/njPRB0OooSWiaMasj8uue/vB9y+E4YgVH6QoJLp32w460jmZEaTxCdEE
u5d5SfRWFPG4jlzZtGuIjuZOQL0gJYuqaicpE2Ws7jBKx1cb5Yobp/pRyJAxDbHqbvUiM0kON5gf
HKFRN37PcmKHgGefsj/V3S2EOwZwQD2M7vdrKvDcMew0Rii2qecAT2B2oTLSEynSfeuBowRrv92A
IOytwCeBwx7j3lZQl7HjTt/mX8UyqzH7lCdquI9o1Q4QAv70lD6sPffskxbjR28H41+I872grsG2
oEGy+7ddRYKn5EYoqMyVbDnSy1/hQRhbPoXrSBi0ClqNtDV1FyBxcQ3yHo1o2OfwXr8y/EXlH75/
dz5cd0yGJRvItl45tyGyFJpKL8kOz5HdQBRx7u5hlaCwjQKvEVvxTqh19mne2CsDoLNA1DTvN9Yy
Ek1adoZ+YK3t2UMphoucYhSkbOu7ehpr5OlOqP9IwbnQyT9dpOFQZiZ9roBkQQLTw4Ixl6/hBpLy
XfjrtHR+pK/MDSOiR2jHvihhLTpS7Lr68FUYQtNhmekr9BkH5GdOj8vqy8ba68pBAXoc6gRsjvwN
0mGXk97Vf235SYgiyP9rkVH0IdK78+Ao66Zzb7ZBIB13T8CQ6OPN7s55ggDUcSiDGgOhglL44ZGY
IwmvsTyFElzVuxyOij7KnktNi3aZ4Nra/jeCjdN9GCQSM6cOKB084GRF6lOn3wv6lc/7VWdzspTS
qkqYxRhB/uV1pxD6tyQcmGIJ+oQWuNV+56w34Fry1YwvkdfsbNXy/tApZQOJkC6yEYsZ4WQOH8XI
tvnPR6Z81w66DRSth99LJfFIkF2+JXcA4e7NS+JQVc6GeLC40pYtMFpgHS9JVHdrOJ6ihyJ8o4Vd
u6OiA3RdJL9DQXArJzemox3HjqPEaO46qLpitFOdeUyhPT+1rOY+kHWYq+LMwVLFoFAKf6X0nVaM
JysAgwZDTEOVCtlXym39JvLtQNDIrJDbJV/8qGSlXmgFAVWBjz6uaYpT8aTQqGNP2B4580EzMSl8
zFYCWElwNZqjkB12qDivJdDozIO9kporMdGr4xydGgB+l2kEjiRbaTh0AOY4YULl/UlAmX67GCa8
a97zA7Is0mWupUbQFETNZgwb37WDHw4Tgjg/U4zDI/uUw/F/3Yuf8sLQZeXFa6bP9VV3+EIzeUH0
AHdDeswxJOChKONxdX9fLztcIuWM89DP2Qb8af5IonVvIv3btIyeXM28pti+0CAN9+Rkv1EcEH0x
bGRUJNV9qJnBeBWX4XI0Ar0lodN9pr1ON1ta5hMGM5BksJFJBH/fJ1JSJFcOcUKqx3q7e1749Uxp
6gD+OXWbGemFk5AjSIaV9+1Kpod/Vr+A7zUmuQXHYYGnovIy1myGskVU5ui1vQk51tudbFW3hq0i
GcLcvz3CtNAHvvdltOw7MVegEAnQcdGd1fXK6fcE39nQlr83iIZRc2Z8cgJ3hEudNgeVc3sEb/3y
IAM6UJQlp6q1tWUkUnHYF345YsDkU82JBLbQB3VjyBGCk5cYwUQejUExGkLlzVTuGb8Msh0SjvQX
zATiTCzOhEmof77PmhWv20asj4BM4XDH2DG7XVwhxdI33H5vlG3ANlWYmyD0oMKl6k1u+pAwk6dZ
VCLEJbyZVJt/0EKAJgkr6Qq/3jx37GMZYY9H0GnRLIjpF15e/amgXUiXphLbU8F8tsESRMEI1Y8g
D9VF8zhU0mAc12q6kYideXF6bNFgQ55B74yy6Yq//eOQnPTzBlUS0B1CB5/vYPIMq9tGjMq/VHK2
ebliyDoF1+T64Wd1i1LEvN/8CJHXgPovgAY5+B0vE4GZRciQkFcJvyleG8vhBfO6VHabeZDXtURs
62BiwUKzbNiMRvC6DVSB0mCl63GSOklDT0psaw/JF3kqTMQVXIKW3BSdrYS+9dyCINjkgHrCPwua
IDJue1uRIyB9UkfkdaT9S8x30Zpn6+/2CavPnGJjPc9Ial1FMTuHU2RIwtMpBWP2bs+bphhUCKUZ
YtZvPbEwxezcondX7WQ63NOHOummV/ks4HDE0CW806rJLLdk5rPT7XugOIk8nYLY+Gzd6SEH2pwd
BkgC6UwhCkb8OztBFmep6TTacCuFuvjYvu4fwsIN0mrtbJnH8KMOJn2LqXFaGgs6+r8hrwzjbonE
Z8IWaFlTYLA+EaqoA0xlo4HBHa7cnxTiB/XPLrHnv86Cnw5fGFt6JOBvrELJa6CzZGTe2LJt1wSn
DFfUdc6wsRpIqeWCLCZTH9ibbSeAXTCq020dNXyTRs4TJHoiEI3lKD6NP6keAKWvD3WcHCxVZU1U
lKtpi8qOiU00SZ13EbB00PhktDo4HcdgDCkGqNeiUK3nI6PtaGxQn76TrZn2ZH3mDyuEW4Jxw8R1
GXiRve6NxaxtRcEfIybu6Ii1XGVxwi/Dm7b6VypsC85PpHoqFlp50j/Qm4uXj5XNhy6k2PChhm9O
P6GJFQNSObhCE4oyNI0vMGQXZ30mR8X7oUZOsuykzXBPuDnf1PrHVn1jl8AeZOEYH+Sr2l6I+C9w
oK6D4EUgKuXnU6y3wIeNXZpjY1C+sbTHOi0kOUx1ERMoYlyxNFmIZRBYJw1xM4cTaOlMJtFgfu2w
YIctoh1ljF7wALljMH9AOYhk7pHAi3eu7OV+OMPhJBrguOP6+BZEOtMo4fgTvoVMP4osmDVNQhRj
53iPqfJxRr2GU4IZ0cZnkY20bU54cImIJIFHxHTBUIB0OQdkYtDkKUbBI407UnidAU0313OaLQiz
juIVpoCsyoOq44hOCu0dL3dQIRS4Y2tE8SSziheen+mDqAcN2zW908daUckXXLon7dvnTIxogw8L
irGWFKpKw5U7MJEWkQkoNgrXx3LtywjVJFujnV/pnVMnY6P2SZpTzf0PsLkeDNjttM1Lm6FCrSg3
cQu41IUHR0VZKXGB6kJprpB2wYW2VYjR6haMiQ1EK3yoSknlxoZabHwIC1Yh58geMBRY5gEgXXIn
F2TCPtJ7ecCUHAYT4x3NIldhF9csOXMXNfk8J0uZ404xpdjmiCr4XakBhes5vn0Pa6/WK6JC8rBk
QfwVjpsKa/C0cTh+Kt0zALgkQ4yyIe6KBeMGc3PZYTv0oC9c80qZyY3Zocte57RDjg7YvcFgE2tY
7SChTDRZVMX+ZAsE4jYg8J5qJUGHG8c0+gMCUOv2DdZdFVRSdC20MEhaiADYtKJe83FODFB3Fvsm
hoa5HlATpZ39ozLJV5J5Ens0c6TO0VKL0jHx99kBobEx0QbBebehS2MQqNIEDRMh8fv7pUiVanyu
GcuZaq2n7R/xk8aUHD8P2NcgifPON3fpskp15fxJzMynIPbWkJzlszZY6aWv/+Czusg2OMHTLR0+
KD/sW3OezRt97vMM7Ns1NtgkEBzF1PveoNn96O9brQ9qrZ8hJd0m2UgJZOm5w86BbUolC/ykPdRf
5e72P97PhDk3rPzMiy6ttzZ6uQkxJumZdtV9QyZOW4WDHzE4sUylOm6OGNlxBP+5tbi43APjnrO+
y52SJwa0W6FJRI9xrtwaXO+WztG11C7H8rodQ07V3iDSi47L2wI6rr5+Ihh5giN4xhYJogC5rTGG
oGOaPaKCCEl18szLArX/uNRF954Or7BG5DYmaVeTFZv99bMMN3TS7KfXmOKqqL+ZSUvuQep4QxXF
GTbNOSEPYrfzXsuK5hOxc++yb3AUxHK/W2MoLDufSXqOvBGzxKgIKA/thGjbAdrF497yJ6S4epvk
krRMieybNSLGhqugoEICyrjSqL7QwHK3K/K+j1/Ddkx/geFkA6B2ZoI3NUb912amhDNWHCjjHseW
dmZbaYE3qJ1i5Y0EOUijLQncsJAvkKdcfKfSBAuuTEJV+di9+rDxbi1lURwwn80KJIQX3t6DuzH2
03Sk5PQe5S4cJmLoqrVq+KH28UqTEeIWy5yUzjPjj+yoZe3WtKXKLI3eOBfXkTJyMZJ69wohHr/O
qQETUZjrNaXuXFGGcoaY9SRN52iiaC63Mlr9V8HBjRGq+DzP371748iKxzCWW0cD9RnnqvNIBQnl
2fbLkyqy8mfi1ibiijvoN01UzHcBVu0jymGa6DyVg8q33mkk1t+ioQMdFjIDZM8plOUAtKLtTjns
VdiHqa3zLNEMy9nDIW0lJpX8DRkfZvOExFa/QOmyoRWYzmXpl+30A1oOAiQ5eRAVboYu6d1cxRFi
KTwcMDFwGhLtBG8OKQgXN8z+pd42KvB+5rI1KHkACdjimJD+QUx2PIERQkH9AOjR/3jCYzpbGVRn
eCPMGL6WCb3bJ+lxDKu7fcKarz238o9bzSno3O6e/NA+thQqee1GogzywdDed4zswN/Hmm1F5zEX
s5+6x0lmAhoo4HgJwVntod2TR6hg3jxQpq9hXzXEVfFICAzsNf/tkeu7pS+n9AjQlb+Gfzie17KN
m5p+J6bd7+PnNSivvMT3M1ExeSyAXm0+8j1qFzkcmaOPfd2yjfakKEaotZtyCSUGJSJTiQ9hwXtt
Wil8Vs7nkod0h/AdMVN16oH/0utfPPkI2OUEDR2CW9XHGAHV8Bpt2VWgx2x2wLY3oE+j81uuZRQ9
/YdY58vY5Uc4o316HOnszoXYbl0Iz/VhTn5OtcNgUi7tvSmWvF3EFfPXjfvSXxadykW2g/5jXk3C
9ns+fSl/ziPPzvoogELTSaVmB0rcHsd4kGs5gh+5auEmvSXK7ZsTeZ7sNvdoz2OHjDzywmF07Lkz
d0+GFb5Pg1fVRavFk6XesgRZ7d069S9p57gDN3V3Gim9q3S72T04g8SLDOBDm2AmNNhYtLbfZbzo
0gPG9ipEvWK3YjLaxxXGurYNQq4O/Lx4XmuYrCKqD6jGZy6UdoDOCceAGaEgSdOYfPiZ6VpxzrLu
nL8eOh0ilQtwTZpZk8eHPReRiQgSOQtWEAtnNqZjLJt6BESP5L7H5CGHDjoiEHN/OuTni48e1zvd
wZk7CnHcbVccRL8Rv+P+BrefDQbQjSOmvkWj1RQUWKPnacYuvKQfzhy10ID0v7uXiHCVMqzmdvLL
wtquqKypoaObEYj2O1tyA8S0haEY+ADPZXvsjX7pnSZM6o3aeLNnZJYoeMc0PmsaAnk4gSctr41L
9pJXVAsH92ocXb6a+rt7NUVMMSQNNV6a43g2RUW8n6iyVfB9FOkWyRf13FzEpt+JXN1pO7ArbZQV
cWn6VEkW2SDdoD/hAQXLikrqu1akTAysT43FS6jPZyFSbmuE5uYTBnNa9wqiO2IwlVSZ8RswaxyD
6NdLiJe+aaW8PDwHdPA0h33NWCQTNlNlSlQvABkwIG4RKeY0TiceObW91fAVdHvKuWw2BdIRw+eY
d3zRFFkbEK7WTZX2JuWimYo6i4ILXi0dxHCagSB41VZSN4tydTWJR6dMr3HinA8tjQ97DVwh8aqr
9Ye3bnjnt7q+0Cqo0olX3pEznd1nAqS2LOFXBnw/ZIQvYwniIFBtzHzaQeNMWn31tQlQEtqbUXPY
xcqhjAz4rso4VWAWHyZV8tfND+GvgoTnURctvwFHWQJbPo1ZKF1KpXN2hawzcCe6XNJJJ+tVb8eT
XMyerXHjQz9gpoAHYsr+4dsRcEpvJr3Tz5mnYgqWK8ve2+lPLUOmaP2iooHyKJ3Cds3p34K14wuF
wnNfTazxCg/+vi8TACzi0I+QHvsp4qXKc4JTMt07qewnVPvJfBHxSf4UZUja/bj3lnM8JoEADJ3J
EXejj/xtjJriuYWhfHa/joQKr3ETWkjZb57mTyYlv9iedqivc3SAXVD1BElJGS+Hc8d1E+IynjQZ
g+gfFR7bUb5h6A0BkuJd1eo1DIlT9JmrPB+2RWkEox8XhHadeXISJfqantHuvuxgnl2EOssEH6vM
FQS/GAW18WtE+/wNKSwsI2ySXfMoshFdY/iD3bglp96mq2knlMyQVb5dt4OIey1fuF5woEYPyT4l
KN1ZjCcuMMbh16wiEKqNS/qQgB3+nQhKvN6W6qF4pdY7PV80XdNK7RimbXBOgvWwX0UZrs13p3IY
nD9KTITQpMgK8J0fVH+FafrkojgU9qJLcSkXuBxVfX15Bm2JkrfyKOymYvqhpOr/6+++sxVHiwGC
Rxqd/E1MhTQXeFUeRX/5MqfacKF/3BR94Mlkp9xt6s+a4TnOfNcWakr/Iu9rL7TMF6czp1QQTe6k
pNB/tD8I+8TOqqn9IWUVXZ9B09sdhw487EJHimU+PVvVWgl+7ciUm7ZPzPtWPg9lXQ0fibQ6X7yW
n/UdEHoUO2kTJkoXJkUYjodkg6uc3iOuY4HXZ/IEbshl8DtcCpZqEbg4uxLZB0g4lzdGUkNu3x9u
dkBJrAnpmkakJIIcjx8BumhojB/TU87X/jtYFc0sD333e0CpysLn3THfH/QF8jGz2copNTUZikdm
5lh5etEd/U+4rBD6n7LJbsAfLLH9OKQheMWS1WvywJZUJpYJc2JGeCDqgt5/dBJOqBr38EC7NeIz
oF7djf/yAZrPH9J1mpSxAZqNjFNE7TUapBkTVKgz3a2aYW0QKB7aTowAmGO+mwasPb4C8/AhKhbc
4TTf/06ff5BUvC+1hPPWRDRvMe9tT+FKG+I3R217hID5xM8BRov4PAq8LEW7IZq+SNpdoeTVYGPw
JJQVjBWXcfy9hMEo7+pYLekZ0V1BlMjldOIZxksr7ueUuPV4J1bNjMx/rAf11px5wnwwAxRZhA2R
LnpYPI1Lwm+CDGSceN9cv5pkV8ItJpdi8j7qRHdXPUIYdVZSMNFdnld/7fgO4bRWLsikmTb8fCQT
SdFA03cHkmIila/oX62oVBxySQmW8bpYTcPITpoG6bqALNkJ5Q2qqCE+6Np7eO3T3LEIfg/9Ns13
gLMxu09Ob33UAevmj3to2En6MsrrXFe2wKHaREe51tJl8/B4xT/Z1SfOHCdGVv+PA5r0pm+469zf
HiI4cjcB+/b2f8gjmGhJkK/Ywl2XfedL0Ab+kxKp6PmdxAeaEL5xAwSFm3+9sghmgJ8NcQ7rQ3rv
EZn/4Dx/ZbgxpbyP5UvoTpT1y0LCIBfeHPDZbx2xrVyTHnEpWY0SzvpVReFFtBYuEs5J0odp9eJU
UELUA/sUh1LOlxXS1Ppox5ES9VeU2KCQacxJtOTuyhvFc+//ECYXSZ0NUtuhD+1CfuYpMoTZztdO
Xpr9ETS4nvCcHQQbJBjXr4Fh7aVyzBMbxQHNde0um0XNAH9KvunzD0EvRp0Mnr8A2BrSJJZ/9HMr
/AzU/4OX2Fgvf/KvuRf0V3+HfoQf/waEW/jwfgtgtbsolM7Mx/oeJLuhJ4c+Tw295e+XUcghY/uS
FswNMxhMOEhBuEDVqfo9ckJbJwFWBahyHHPeGQJ29cy9WkFM/aFSLbnQ1y+Qq9+n1ILTKTkP9UkK
VE5qcFER5n25vgV3O3WgjwvDiw1NNpfEGWzVgXA7kDRuI8AUEizl+Q8ec5ZdeVOzUiwcH0O5zBnH
rwKQ/K8//Mhg94lZ9nGIPXIBw21BbAoNXwEoTHtTUqJ5jxRkS72kthB1oxLwdIo2uNDoKAOW07/q
dxAl79ugrHnMlsq1K1fMeJO0TcX2AqKYps66vzgz/RdhXzlTyPbOD+e+x7aMApwhSAOl7k12ULgh
NRAVkjSN5G04AC5xs3pvJqOuhoqUltvdQeaNoDtBGW+U1QfcYyDh5guKr70eMrC/MwGUOnHnrgA+
2S9coZVM7KAD2xmDRoUMquKStfbehG5WWf33J9aqYwpZyjYI8z4EMIyW2c6T9FCtF5at00tjopUH
JXdzITBe6yQLIu0OKuCgmLFmOXpA9nAJG7XL0Y7VOwmWuGML5LvcnVCLmZisxIyfIFqkO+/t/xuc
hJ30EQMOoOw2ZQK6Pf6cvxLp1jpUDRNbQhijPtexXjKFG7rxFAJdDlga9XB5QYzVydlkKUWT6XFZ
hhJurMTLeuoLCm7YTiSxlB+PcnQ2nKK824GuZbcih3DgU3C5g8u/mvIgauSRRyrpemnkVlsZmWCa
e/iR/pw3nBjdc+jaLqGwTH8asfB89cyFs7+I2MfXc682NxJ+OaALj5Utg6lVimcO8aw1reDo31ep
GkHqMa2JlQ6r0YpzMM3AP2a0qR0D4GFtZqZVEvrnLa8Hkrli6S4IPRf5TPof2Uf27s5DXzoaTJz9
8eNqGBXvnvC5EJxIwd8KTrb0ZVnQxuscBAL0bi0lDrEtmM+ikebq613HxCmXvoFBCBDwZAa95PQH
vrLVtc9+ByBAv2uo7DmADshke+Jl/lGqAexgAsIqmZ4yiVCVt/gP2wx82LI3MdGBQuB3PSxC4sqq
gDL52/7qW+A7V4jxZLxJCYFUWY/vJqgsoqBD7S+Px36aLWEcOT2ekseT/jI/sVdTa4EqmPYNUncO
4w2M4d9g0unSHSEI1NCjYyNIB89sUHRfdn6CE7dTDYpUGtOswldMFAbSObniJxhgGlT9D+2/Kcf6
WkfWitk0UI7oNngsq0fJDZwhh7OfCYt7BPbsd00aASbrp94hBW4K0dEg6VWbnEFiiw3TkA+F5h6K
mOFzjMzsmqCYY2eyTbGNG+2bG2axAlltialfkFJ4nQ8UMQRLud0z+URE6kgoyonD8hFe/9AIpdGn
YLkf40fbJ87DYDeaaSB1kAnzsxRNWVTmsJHixprfrndtsscjMwuBOp4vj5I/AxUgYK08xpNwXglQ
CFuiUngMVV8nn7evsnpFfLROuCUJc05sJKTHYB3AS9gqgCW6R0H/LZ+nKU+datFps1vUlZG7EAZY
HYrRUioSAV8AAU6XE3Y3zahVtYwjrgISHeDsbXcIy6qeddZqjdGsW61oyNfjpVXIiXQEUpfmVWpq
UxRUBvN5DEDj8kvqk6y7x2Ac01AOm5dlSoTVhsYxRdn6r2gEK8i1FZlrk4cNk5aT9IAo+BwD01t/
9IhfvAKTpYY8QMp0c7Uqg2qOjVhN5cqkxjXKqVxf5H+MdRQYI7BDLpWomKkQlsKwe7ikojHQkcRm
DnLzMmaNiHFu4NcZXeCVt/tbTwHTlXoBFZOcLtfn0681qOfuYFcOgqVmmWcWMjGCMzBsNiilnysp
7kOIttzd8I7HTwo6S+varzev09ZlKwD1HqIshaqo7x+fEdmTdanJAWwdvK9Sp/hoo/t9Ndbsd+ZK
MNe3d50UFUmQ7FiZAGwpElH5HHMGQ7FeAsKyStjddWrYxivvwMyp9yfcUZMWKOQGcnwT8na3QeMh
huxB+oY+7Wf+2shuTZhpURtMukcQOdpJPgVcsgxfvHSVbMSrOQ8h6bUvIInuW05OnMhTvjil+aQs
ZpR7WKwRhWhsnii72HWv807hcOZkUGansyDlLmxK+IwQvPgEgVDMOTbV2+ATHs031Wntzh82q7yn
WhmOkrwrmPWX+zx8xGDuHmk3BgV5zu4cgznRUlIG1t+l37QdYqjaovA5MW70lXFQRwnjrU288WqS
Qn8y1dlHkzlrD977Rwmqu2JStPBI4lqtXc1GA0TgiecXsaO2pfBVOZt8vgtLlU5ieDbaWhlPVO3u
5j6fULDkrKLX0xNZ0of93INGPrs+2lNeuAyZlonPh4mmuczU43qc81NlQYDwkUkFDKz1lmBj8Eyh
B6vagiocdRIVO2x+4x3JDdDkFHinDRmHNP+6jDiXIvvMqvm40l1rFkz3zLD5SK/eaQANgKjDtQCd
wud8ojzziHrzK+ctPWYlyeCHToYStoXQwFNbHrjd8W+osWGIiI+CzXEB/d3TYtbjsgmYH+TQbcYP
05qSJxWzVwSCbxYLAjpV9KacM3MyQJTwcZ6ODu12OpGYfP/AnSNyQQPp5xnh22RbHHxXKK6W6V9O
y+0Zx1T2Zmuok5C53U+9aJU8nOY33f+ERauPGWdRpPBQLaOgkn46QBlQiDwlFMZvkMXL6CuBLf5P
kWFK34sukmSBeG1lqUAYZrp+EGFnXj0qzw5Qvd55s3IaqylJrVVY7wrsB9/CDI+Y4kWovvUbqPKe
9HV1ahaRBsevqMqVYVGTxjDGYLL0lRO1OfTNhC+CK56j37H8ZhaKUeQcN4iLzGD5DvV0lAMs5bQR
iM4Ir355MCqQaBwUz3V9Bnr7ByGaIPaY5L+ChrGs0vqR9Af7uQLHWK8B3kzZwsJiC3KCxWtC8ab5
bd+Q/T/esXbwW7KDUm1lWr+GmmQtwu2TCPnxA6H3D7j4qj7IiUmU0tO7uiw789rIHolbBCsmMkVZ
Z6C7RbTxE5o+s5PdcIZDtlLa0WeDIUkZpqH6mavghsw0bx7fCtHwX8q+8THcWIjFOP5fimY87LzW
/wVw9VJ+FUZWpcsNj5Cg4NTwP/mz6Y2pG5z6g1BC1EKqpo2qKGwCc7hKA1FTE725hVksRKBkr/yF
00L/UJpObpYJZ7RCuBaW/+HrBzlZBFtzjbMn6GM5FQMqr2QoAfAMVBANLQeHY75vaLCbpbFsnNQS
wEiVWc6s5F526vqtri5jIDA9OgpISzgL7Ar+vqarPDREyWF2YGuNljbignkjlmEL74HSoMVgSy6j
oCOYT0ZpCxcprrulYUBT5mZl05uAiGuUMidbmBoNuqNq1YZPYcMx+tY+qG55o/J5YGmK9rOfbalV
nKJonQHbhN9qF/GDI5DckZoLUp0g0wiJNVr47MROgsy0AvFNHalwi9LgKSqgBq4pUtqShRJMFv1/
YRteepQLimj8BUxy0wGvgt5cLw3XaXeIaKmdFIjZevaLaPAJ5BYEFWBsZ20Stjv7/HVAdtTkq3Z1
QwSHJwjovdmgFd7OJZxVT73ihWhx9OAwOy04Fzo9y+P3kpyzwfWJItuDCCqPNpCf5SOg3uL5s+nk
f528oojky65190lLQx2EDLgB0oWUgfC0YT3wKL/aY2jF3dbUo2XZZJg2ptaLKxfWtOxSHl8ADoC6
9H7U2go6CtttGnEU/abin/Zbzl2LchXxOJadOPm/hpYZDl70IdEf1Qv7OutUVxeGZRQYNfUSrp8V
7V5qZ11OQbGk6P0jwyl7Xd30O1M7Tt4XXRZ5yeWjN7j4kRu8ue1hh3fEfPwvL5PNRvZKiRhfDAxo
203nqrN1VH9BCr62oFH8EZVBB1ia0exG7o5Qxnxm/DFhuzC3rcGIvP5ei1IUkscGsnz6mlhHtGJ7
D2sHMrz6/7Dqiu/bnexMbX5IWmnNuepukIsXO12e2dDxbQ18CrLpGAc+mXrxcCqra2m/zXIvul0b
oBL1ZYC1QW82T0/RvHWtA+S35YdFgpQKHWZZMEgg7ias1Izl4pEeSzPr64HfKNyYYtRAPeLPYoJJ
6ePd3eFFx8h1sYGJbhSxOu7RM2UYb6RlHmxG4fbeAc2v736sO84hvwVi36p51xtm445AiIIr1GRH
FRyFcjphMgwEbTVQB/p9akG0WFCO0dMmjMjGE7ESoS3AIuwkQFigw6vCGzMn7qtwaEkUsst1isd/
sZWcCVtQr+e+1lM+L3KrVy9tWLk16XvDvQJ9gi5pZBaAaKAH8zzkyau0sEwd/6G5OWgOzgMBGoMA
dkZCoyV/Nk6uyDlob+3Ti++/YXslB3/KM5qpn5FNjKGXy0Odakahj8P3M1LN0HiWEqdwNuZ1/7jT
GuJdESnT+PLHv4XjjWAE0/VWYxi1v/MYwSoODD4RA56E8k9WmxLouHt/JUViBydrQaWABs+X1xKD
Z4APPMJDgcVjHPowpUD1zz/KQtmtxZaebrlUH1/qwuD6a/cVxrSQOdajMisUdkSjV+1p03ywOMPg
noORyabPrhfqGVkJ2Y2j5JZQfVZqESA7ITDSB10bU0zn1v8mmLDrHh718q5z6n+PFqfTL/sVtbCP
OwCutez321BFjezhogcvACXSZe/AukuBUTFQrWRUmS8W6euK6n3MOD9U+nRzNahzCZTQCLRkz+Cj
fTPBKHWtfl5/2yOZVaxmbsVDBbPqbs6uwZob4ByQ25dNwhcUh/fOB7q3Msr6HsuGYGwTNZNG9+g4
pncjrIe1lk8vNtl5rrG+o2vsuRo1Rs1QOFDsy3VSnpbeBfHL3mGRjoIXSa/nxjkZNIplwy5DNnB5
GD/4Sp/IYv3I0YCnPc8/hmvAqUhYFgtg5CIwPmYwKZmdxHZUeybqyufnd4zlo2psb+qvZqURl9r6
5X62h0kCo2vLV9+WsBmslmI/1jkYPsENaAHzD+TgNxmzTHk26293EqWTxiV9xITZmoUgsr3dlnFn
UXBj8pSwcQDMH4mxPjTY7EgNTVehdTDu/Eozxxm2w/ydCelr70Rnut2WtQeSchcKs1rC0UDjHBww
v3Dibvf3WgfFjCXpTDP7jNdpoyPij7iCMv81mLzprqJgTDoc2NaE6MDg/XEle7MfdG7gmHpwGfOp
euJ1Hp5MiqRV+zjUfgT6/S7crEeOnxue6SKGSBZilF5qd7yDP1XnZsDx+TNUDdgrfi1Fb9pW2cC7
ldYDPYsS5GipUmlcC2TCKO66LtsgQPL1OlNOXcLLipISJS1l/DpTmHSGbwziDRZLHxPx1lidHaBf
XrVrhB/CuyGQZ+AEq1H6GojLYasG2Vl3rAkL4yqk/HHKcYaItpGCT1+0F2icCkOsHTLrfyxIWZgf
u+DQv0eSFEMP7jO4qtTiVxx5qEm6Cne91LuZ9tv/ep+SMiy+YadM+2/INzvh/4yUqQvpdf27DN2e
qt1uouukOCrdTDyPeNJ/l8YjMhK6ve3AReVi31ZiLJyLkrw1VShJFaZpGLxnFa54ic60eQuaBjlp
iVTdoQxSBf5LGhrDo2teVcStdiqUoqOHb7Ykvdqw+SSzuit1NzHdaTHIkc3jejok9FjIvfSnzZPs
21H+ykFjnDttXAUzMNKfxjcG/NvKDUkl7vYX1ya6eMzbivXgfrlGEvKI+wEhhww2rGFzf6hsP0b/
4Fig6NsmYOTCey68NyHL4jSHyfSEEtDero3v89PLR15wZrXti9mH3Xrs2WYiMqFx/eYkvFZHr09u
us8795ZI9RyE2Mstf5W3yoYW9rH3l9A7lNrhhTn7ExihUnzQQmyn8q2unZvkSQ3ANImFxLX1BTW6
pqc1RYezfZQpZ9mCwx6ZGmZX9AxKf7SjjQmybqNOv5iCEAdYyzkX5aRpm7ftKsehBXiB700WD6du
fdxd/DqCJKdBAbvQVA/i2QNZwffGnC9kudsjSFm1bXVwySdK1VXg9wihgjvxmsTkEHJIu8rCXigb
Go/3dGsWUScn/AMEHIJm3P9ZWe4CAgDthS7I2M361i4pSmB7Ty0MnUJatWiZYpmvsre1WM5LNzRI
qdEnsabFo9F33hIapBD3U/KA8xkSa0DXADKkvyYqJZxEIqA2BT5pZS/qzblutO6nU2lx6VWVfl3G
4cLmpNWvRXKKR8QCF1DW6OsnqlHtbfVOe35o5aysXA2NCwOGvtlptrr2mYttNyOa6ZjRxJI2t8qt
4Os+w0cW4xbDGKLZk5bGcWi2Uhk99CUZnPE9hXlbBVwhEI4TYsOp3PDpwIyoSea8WeJmAjTHYh8s
5AqHvdQT2Nhf/MvRDK7lh4wSO2DcFM8wqIb66MFR1GsGCtJY386KEBkx5huSx6cDBNWMhCuzcJug
mk02Hw9ToFzuDUu/M5rldXd1nNMQPtu/ZMXSXUsTb0VIyr0RCPYp0m1XiB5CwEpmcxTqCD68NWqh
gsrv+n9wrljStHxO04/QvjHDZWe33RnTzjRHSSUGnVZrPvleKxlrjFRaOtC/bshHI1YsCERSDDqe
VF2K5lD6U7JDvOZXDkaruu4OvmxML8p+EsbAIPPW/Oq1llMF0dEEQR9J77ElYeGTvK0thMnShz7R
UnPTqVKjmvXS/SmQsIjt+rE8EaWVysvQdGIORNc7DXnEObq/C1lZja8HK9EeIkXT21vrgKgLqLBS
FNJd8MYKZDYqqwGwXr8azGz97pr0xJYym/6Fm6IDlh9VUZOpR2KldLQCq/i+bJQ8D6qWXtINBEla
cxF/YiunT28OagH1OsyB9GB85gMIlqXmkTXRWeBaoIfb/Or4r03bNUsmlZiUH8Bj/jyWYnbi2zDm
lT+FKxTxtHvZ20cYgy3Jc1DYCT9rQmchmh1l8jnGavFx25EcTRadnWsYQ+6qw5BRNx3WMZcXIoCU
hS8fTaAwnz+QGKBkX4nWhJrHtAtWoyiZ6/FPSdnQSEagIOawCJinLl3Ay0DzehIGaO185N16vjAn
/BQrZNPPVoqwb9BuOd4RnFZL4cRGxrN/k8eQ1AlPMunj23LygSr6ijw9t2Z20Q/knZUss118F9Ke
St1vL5LRgn6HU5SAEoclyL2Uuzv2wOHVSCI6EuHUmRV2s0wgqOn39UD/D6yIRcFK7gDdjIQo5VMM
F4UtXEG9pk/HxWZB8/eAbhZjdpUbxNzVlnDQWtQzEEFYHAWNwi7JVpAWlaYOzP9XbWLnueQ3Egas
UJRKh+LhWIeUQqCKJEZd5j/vuXMhdfr7iuhHgpbiaM99ggm2nBCjBkQCRWv4dlpujY/ftjws6l7h
SVAHz0PmRscYPdp2wFCGJyu3OA6EHYWjhHYlYlHQOwi4ezX+gHbur9xzYVA45D8bsuq/nilaXVZY
sTG8X9UEdA9GbpvyaEXmlw3GbLjtuwtqad+STLiyxo1Z4GbGla6APKay6EhZMA4kgxYB8kPScUlz
xWyxS4xCPshWNrlc/DaXSDRfKEl5ukMs6Cz2WxI1AAaPl20hNOdgKizsUQiX/CZ5xu0NfX6vAssf
E68Ue1T8afipv5UBx1fP6MfgaAD0kRUh6jXecwjNuQV2vyfAFwiGhKiUPY0fodP6UZIHtnwpZG//
21VC4/Td4mrRXzThcsw/zqI7Qgb/GFXTzVF0mAFz9z3gY8/cC/oc3iPEflFP+StqfUImLzAzCu8R
NdnlnaDqm1Ozb/xvpROI2aFwvssGsY9BE415F+a6ktfoX0sTY8pAkfgO0wo2+M0YDfLxh0Hiuwuw
K7kR0o+CpTYllxr841cCOxGlNCspMcsTEUZmEh+eJv/zW/61bZVw1wUGFG1zoXMnWRTXYaDh0Shm
t0FuYROX+Qwvm3Ufuul/JOchaQNBp674lNEy+UiQJQsdM4L5Y7N8MolhQ4FRmQJDJ3XB/8SmwvGJ
+J6eE1mP64dnLS9miL7QTCP/X03etxNqEvW1IY60eR1VtY/AF1/v5HvLafPH9XKLn2FDJpCnDsDP
B/Iwm0jQcn39WgCApg9nqyUdJjkYi7wh0yThuQLRreYtTkamjlAZRoaO5TEaeIFUlrwavmGLS6bD
E/esm/LIFPBY3Tk7jX3/vmnmQ20mUfyHZ6CXDQx9IfTml8tqjuv4DRGv4N7kN8Oj9I+piCauPgdD
svE2cjsf4SGCKNGnhOpZrDEDJROiT+HG+ZdiPV7/ce7VOoSw7iY5HdW6fTvCitMRY/FHrWMMmU1u
BvZyXzMA5UFxoJnZ9KggRYn9cF/uHYafrSSj4lmfo+xgZvnLjEWJZQbR84wpUwzo6iXN59MYoS/t
qso9YPKstHLXh8t5uXa9KxOJfuT/sDavETzhDF03NeCWjtxpfKJUlTCjiN/NUvVJGPvC3xCD2Efi
4f0BEd02/MZQC4sQqPT8PC/2+XE0lDtUto67ydfFg5FlbOFfYDRICg/XQuKKy335XgzA3NX7YoOX
UJKS9EcreIfI3Y4hqxxR5bvmeX9bX/OCpwFhPXMxRC+ZLwx3GwPnk94QAESsI7sTmKmFsj6mjiv1
tDSKfAZDQFjHlpJ0bZPhALX94jqGnjM6GDBI0hLp2lJP1zDPd25MEhVS+QnVdhwUm3r/1UFYqic7
2tMbsplD8CMGOkNlPECCVHxf0JAJVZRpRn3BgJztg9fpQ8vnKaYyr1sqt6lLPn4wrdubrxDR+4bT
DO4FGAOTiX2mT7bfoXzU5RXCG9elt0tP1VICeoX2jYteEKqH4B//yltat/bcqlMVClh+e5yWJ6T7
m7TdEwvs6ZzK2Zzb+vlTnFK0jnJvApLcCWnHPt4rIWAo1BNVsnAjEWa4CayJ5HrjmMwKERX+AJ94
E3S9WSfszB5B+zL5v6kGpBFY7A4kxiTYzzrymVDPmXcC0lXJUfgRXf/2L0JcNagMJ52fFsEWrwHH
yA6CWhMBA4hWvy+/WgZJep8x8lWaw8OABMnbJOHjI28vMnKURy/OlnkWGqsTbMQCSET09iFTaFIW
ceWyUtiewtQmHBUBJdh35gGWpFsRE9PTOabvnMR2Zafa+SSweqj5ciuTHKphsnx/yv6D7aRNHQ3N
oOdwS8XyVL/JLAFx4//YexqIlmcU3BUSR5FEdy/5vi+nJ6E6o57eqvon66vjt8k5jvmYLfmu5LOR
F4uhE/j3M6ax/U7ZDPJvKglfp9z2tey79iNCaOulKs9vNohAqwV/XhE9dEyf8gKKOFltCAfUudt1
qtoFl2FY06yEVjfMztS2tGTHbbJEYWSeBx6261HPcB3jmizryZNzsug5sI+GmBprHDBP+RufF2of
9R/ghUqvwF9jtsG97lIhO0tzVflwk40ejFyZPFJGWPzrAIKhf4ue8rZK+PiL/GVtlAGjFHCjKDd2
9DIncw/V4s2G3U2jtcOHUegpNPs9ur2nVBNPjTr2+e2uwsxUHlwwuagDLsieE0ilS+wp7O7K/J5B
rq8vzagbNJx76/ReUMk1mj1GeBDV6WP4mImj+kBseRaLD642t0TI3kA/EAz6TG90ZhmYgIQPMi7I
tGddCSls5jGK5aTFOlO2GKiOmF1Bjmwm6wkEU7KlRSFX3dq0W2BSi3W/lYvUPDPq/jxmdB1SuVgR
kh92bRjuqhQIZ+Bgff52vK4ej6Nof8nsVhTAczQMFFDsCljFQi8Gdooo3an3Lgqq3DVssLlWyodf
Lp8PJNGY7MwFMkRDzYrPF4WjLhYy1715HyG40L7LNBUB7TapNjFRCi1YD8ZVngGV9guH3u0Qiryu
z+gB17dBaSr0dOKxMmI1KQcBWcnreDmi5r1XxYJUmMQNxXqPDUHh1g7y+UbCVrQ1O2pgf9D8nZMX
1W/z30DnfeUXVBsp8Nq2yux3fI7eU22qNYsMF2QpyUCykxS77YmJhSAxT+vgoOkYANM2Qmian6Qt
M9FLfoRb9Ii1+50BTquD9zURtYMler/iWCW6wGxd1UgIeTx+wEdHjKxGbfSQ+zYDrqGcCcYZM6hG
1DJyefayiySDyGCCzt6e8IzteK9PkTkcayft9vDa/Na63BMpkFCk1AC93UrJdNKKJ7W9BnnTAK2f
xpRJH1If4SnPCZps8FABYCiXpaBQXO29Ik+dwfpfpHHPo3+Hj3LYLOKAhL5+nFdNMDmh8D+zVs9t
yYPHmiuavnGP6QY6WOM18Z7foX7/kPi6dnZrG8m3jdhKkXe4A5YscNnU+SxR6elu0/6ZW6SOw4KH
ar3d1YbyrWoXbYRVJ1dpwOxCmbz+00Se6BK9NRvuS6WkO1Koz2619uJI8lHsXQvC1J91J4lkd0Vk
zq2taAD3WmsUO/IV9j1atr7Ba48WF0BTEE+KtNUcbzJrBz/xM85cPYFl3PrLFYjM6SfzvFbNSPWN
eBC9mdziMFUxQ41mUnNk/Hcl0Q/nxi7IyALdOTqcWIcFDgg1GJmrVi61QCyYVOBUmgtwOvcJxGV8
J7VVjz0zmv4bNEHJ0cFZ00WBdVK9Vt4EWZYkja0uFBjRb/9t9TaX0zIwYS5BRcqR/qbTfeG8PehI
O75fG6vPZ2W4Ek83MeGwt700kj4RurqnW5XzqDjzqCkdZg8NJkNpVBRxgtoXsoBMB3EJJrjLFTVj
H2S9rkQpywfRn92YToSocoxjC0x/kSsGYwUmFm3/UBSRtlgo/Bzepn+dUaKtl7Wn4IP5X8Q8xB0F
UI4Art8Jp66466cPQqQSBu1JBjfoA/xs9YL239wP+8raiDETY7UVM22S50lBSa13hLMhfMu/Dgt5
SlyLAZTf3wpZChtNuJt2BPure2ENx/MqCXuiefjSkvwhZcYauZK0q5miwudGOt7EnBDuAMjlu7U0
HKVrtnM14r9lWgn41bYQz7x+T3irb4fRXQ3vqgssQ3acvMEFmpN+/VBMtEroiiEp6Tk53nnGYZ8S
X+LGgnnLgTR/SYT+UwCQe7E1ZBSZN8zIF1E0AW5y9PvHGBX+wddLM86nw0pIaJ8ee8yIAQpnXejw
0Tl6aZ6YBw7qhsfZf3LOV+UDST38U2G3WdWx4rwcKSe6Pt+fxl7pJuFMRcScueEhPGJ8xZ0QwXuf
WJdMDuMV4nrMNI33t2rNGV5Z0pwKhW/G6AfSI+mAV+p+WfmgNeeSyulmic/cDRd6gR+q6qAV9lxO
yvQRl9syT9vi+ONRV2k4zR+YdYym0LKLsNGRlQvHeH71zk2GswHVr2wbRFdJIQ78V7VMyQceDNF0
e/PffDoPWyrB6+CQRTQMkDyDiNpZcQT2gEzC2cZ9IjL6F8QlyO5uIVkHxDwapJluAQ7DqjPbvrtZ
dq9Cd7pmihtdLye1evDwPa2NNFahA/dm231Y2Kw3kVCwWxL5X7GgV4NPnO80ud+5e3ZYcgjP2Stf
8GRrncEQl3Rbn4KrEqU8qCXuMKPp299vu8SiwVn6v8LBG+LTFf5hrE/DY4P+qoUQ8n9UJVCtq97x
JnrcWFE4tbycZBxPLxlDB/nu+4GuXngBogWweeNPK3tKEmcNebvIRKgXApHzqxFLbErV3oZLJ1PD
D73D4sNrfGFLSd9/47sbWh9R+oZNC94v4BZNwlW40cvf3Zrg80hCGjn1v6c2d/sIp9So6UAILGGr
0JQf90DQMvMgqrZvGPNerLJr+sZnXNsxkOyKKAPiAHwOUJxwI+aNJfNwS2lZ6aLsV+MZuzfNhPwj
i4CkkD0QxM16PyWBIbaJ2djYuEzC4ZrQM8VD83UGkc3XnRwQnnOTXSSe+eXpHBP0VCt85RnY9Hzv
HltzY2+4enxYEMNakPe2xNQEmVX2fvo5t0l5ne9uR0bQAagEewycBCaaUt0n68Zk7Lns8vItzT7e
kAfoYiTa3C94aG4fP0fdF1ZKYJ2d1Bsbu9aOIjIl139yUnnSvO2tZ7m0JDszP/lkWItU7YkoK21e
9kUzPm7eF4EdiitSYcPbn9NMSoKYB8tCs2Th6jB47sLyDO/wFPfUhVi8BMOVlIuhWy9BmVPlI4UJ
1QG1ZDW8Mt70xJ+R3bkc7sy31gPDYzps5fVh1Q2wSZes9CTShzwmXO0+e2s+KcENURnASz9Hf28n
3tp0xuuRIy3G4qEvic35fdtswN5dn9FY+GgzQ9B6+9xtaYo1pQgo8G86wKqGQb83kgFe79gOAobx
aScoYnhb42IzK7u4GD04mUtxRXe8PFG0sTj7HUybpQBidgl0ITEfzdrgTCVdTe21m2Tt3fgNgOkF
RGzQkO0diSLvniJItAf+TBvdU74QBWkLdsFIr3UX0n5QaU5e6cCxjz5BJZKOyyJsz178VnqDBVkv
ciEeLx+dYkL3+CTGcXwCw4D1Lg8YOynU73DjpIIHS8fwSnIfngMMlDBpPcft9xPtW64OU5GlOlOQ
Le1G1xeDD0vfprWt4UGk6eYFAUmpl97CxMBFHdj+kJUOWEvC2RXyGZzKRgAfYMFt68FNL7rsm9QY
OKjIo6FKiwC8BXrBYXCCaWmb7H5GVbNXpQGWxU0NvvihGQaXMqysgN1zT8FMBsm9/r3MFCW7IMPs
pFgXOzyv6tK3HzQLFMfEvtdFbAaHnEEJnRFZVMQCNJnMwpd+08UHGkLaOB2zzDVF3hT5XF6VxEBR
uj0fO0lPxYUzZQyrc1QSBwjfbt6Z265OM+bglGeAHVw2tFLLbxSolaR2NiBfVf6/ZEUr756lcyfp
UCIUSuzVzNnSkV0SC7N3mG6SpB5sFTZcCcYwyyauAUeWWTHGMgFiVgvZsD6SqcfAdS7cYeaH+Pqn
uKidArO4bKYO+eH3i8d7NhZ/gFggiJZK7sKt+ZNbMK6N1c2+fBXGoaI7F5Xkx/0wOd9pwduKCw6n
3rkW4Tgu+ywjZk/AQynIcOB/k7H0dPRae+A9rGxLfNyUCmCV9tCTX2MVmuzvF15rqzfxXmtZsZIL
LRKGVEiQy9lHiXhYQeX1IPw2Py1yXWuUXHluoWZAwNOaLxVzJ3HrZghC5O8+vIS3RZ6gLraeDIJC
TOYfJ0AL0QlilvkrUrcBw8GG3X1t5Q+gpY6elIvE9eZAq1mikfl4GoRLBcNr0BTXJRkdUyOK24Ak
Q8d/hdBfAQM6nNqa+ZRMFxm/B7uuEFdwGUOe93HQ/D6SdcNcWDu1xZ0qDMc7mReA+gayGunMO+tm
f3YgFWOPNiVWg0kzK5GyXaib0Ri7HW/lIMj3jsEyllhkFuyLI9D9wJacApPwo/IzGzV9OXn19rNB
xusR9NshUK+/T8h/XKE/Z39Lbrxuj+5S2Dp1qgnlxUbS6SXrRRxV8bxu8HM1Q/7SEIIdqa2E+LMV
prJcu6GKzA8PWo0FI8teZ+BI6s6FWY8L/4WpWOolUNZTszGUDQExpndiafxW7nyuSn9AFnnqTKCW
XytSN+AJMQsSMIONRd4Tfdk1TcDH+oKgyY6CF2NzYYQIMYYFsaULRHbTNtgG/Y5CGH5+h9XFEvv3
tqJsIkAuRUBI+d8tAMb1XoewzQ7FVJvfhq6TKWQKDBo7Xo9R2cQ2h4c07bl7plm0KiL65/9XdzPc
rZ8YvDCxhti4a2tUXz/cIDHatsoLCMPwYsqw5PznW5wpceewK+H62S5MlNVLxnd8pLWmyNAfc7B0
ePx9GV2bNpiWke1un5TSOCmj0HVlMLVHln1TF3CQ3IiYRriY2L43yB6eLUjwvGVMjFxT3sSgSoDC
mhsJNCLgdJbZfp4trKZd7meSgHoCznPppH7mVPveuRW/K6FPA6eJ9SoKORTbsJBHU8N5KVOIJG6z
GxcT0lg2imJmfkCXlbYq8zCVOw+mi5v4yEHmArfc6SDWvOS9M2JPKeAYZ7OMTq9uF0qsHOqnD3kd
YXdTgXeu2lsxNdobuRtP/4FVspLpsPtbxmmbyU823JlOL31+1nyeFxyFWaT69H/ntwW5myQbfARo
25cvHpurQUHfc1oUbmXCgF4ML0NxgTQdKAKflmRFM1jkYbH6Uqvf5st8TSVwsmPLjJ15KgPCn1Pw
+6t5q7MHOd4sXXCxKP1cDV/SayUfaFsB08o+3WoNiyPbpqA9/aU6Kpjj8menKfwDSSl7lOwG04LA
o5e6P6jp4y6UQMCPaG9MOnkWVMX41r+C1cpjjzGzdeKoqPHnKI7wsQIYYuI2I8pzbL0FSHJhL3NL
cAE2WevqjGU/5zL+56Xc7TDSPebGHi36HEzhciTRTZ+cMsej+TOL9Y6JPX3sWwPDEtalQY15S6Z5
NmrfCJQgNEVfw+SnQpJ6lTmj6yhZWTkzs1mFAZu3f5MYf+amJkRP9YnDelczfD+PDqa5OhriS4Ed
uQdy5kgyIU/Etzd7KuwcyvLJVfnMU2ncUgfRZClRK/YzVT2v2j62+eYnQy5ho1dFXjpZp3RceEyc
6RQXU6S3uSfn2LbGvHp0P2bJrQjl1fDvZExucaZirihuHkQcjfkbeB1teCXqb5jmTiNGC3Qk57U4
aop4HPuHZAVUL0EQ2FahzOf3Y5ADO5V7BhU08fr67SY9P7xnInoNrJ5fDqLkUukwbzUo741diHD5
jEeHg0BzYEOQqLA3FU36RE33EMPSF8jHgkol0SLllJXYsVfYJSK+bEUCoLQWtWQp+dgEKjXKuwlV
wQsfwn3KyCxiKpec3f20BJWhUOPvSJuE6PYUt/2fQCWEDkMvSkeQftp3CZRbRGjPtY4kqUN1ZCeH
Eca6WtaMNDGF3fk6nL5uMxOQfahWVABqvj0cj6xpex+aG+zMGV8EVkcGEdH5SbvnoiCgEhohpPab
jJKIz5+AJ4OHOI25HqsJxgq5qIOlarIEwEDkfx9ma33++k2m6zKFwtmUDS+oqbgsLxWmAUBH7Wwa
oyB3DbtNoky3IzdX6uZiCqhD1sCNN8l5+JVpooxXPvql5T7qn6tqtAd3jhxltx6/xeFZQXLo/9NW
XUsOuvMAqPMt/kv+mfggVir+agn8HAEYc23fvmG/1HZBfh3V6Nk1Iz8h02Qk6BGc+WBmAlzmgDPw
DGLcwtDfAnmLzzwJaHAIw89pAX6S6rh6qeQo1xuO/jyx3PTCD4XQHCl24ubggNOj/0IcHKAsj+M8
8JKnELmAh0L9bDDfaC8XVTBwt84aJrwiLRLuRAKyJ03da7rTcBF0+y8+b0Ls/kfVYxVz49EVYoOH
mjoQ/tpUQugP4ZQD5/Pko07C7aNEuRe/Ll+DnUheXJ0UvkkSve+1CGfy0gwr88wIDJ6wGqZa/F0c
YlW03AnDRYzoWXO3W9QyoufFODvmP3e6s/35gyPu9dCrXFx73GDTePbPUvyor65OCv8FRhHpWKlT
tYmhZh8pTQi0MEYFPLeIG5O2zoAuaLd2zHrd9WaKgZ5lF0s+GK5goSW2n1h4VWj3yZoY4Yc38nkl
8+t1S6iXz2hT0PRqQXpbiTTzy4nBfZNSeyzMGw3aMp062Q1aaS8dwxiIVh8scD4zK+H8DEKAdoSA
N2vJ+uJu/O+tmAcsqbsbxHjPPHDh29fyA+I1twPBDlbsqAA2fWtriAgsen/A+4WdQ918OdQBEx41
xRzefXYnqKSHyWKlYruDE56jv8sXJ1Z8midw0rvM8bOTLDnt1mfHysO97WJd5cF3xlfFMzft6x+9
IJGO5fNamxWhHIrUzj78ikO3KHrMm71YkkC8Vk4Jh0YJjYn4A8vpElIY6dlTSCyPjRn1xtSlEG1T
/yXEIn7P9oUO0B5QIunUgSzqWDFnMZubMVUwq7YuYg/gGRtiGnXBBA9n9plffAlw0tLq+1KPih9T
c3KbzZ98Fp7L6K/mo7Gjkq4oeo3TonA+kWFAvq1of9H+CQh8KWrkBETD3lR1pwlSJk1Ky8zs9tY6
zN+vBh6MNL2MYUWAM5jAWGCn4VM1XbjSqmYn78tW7bcsQQhttNCaTEuLeBmtqc9nLMqodKyNUoGF
TG0Is6lX/YHhyoa7xiUEZlTQQpoaoKkULYvhHdWPM8HCwxst+6YSuN0dtWaKUOcCDDVzuGFNTkLM
u+RGly17ljyyDFXpwq1SQPkvCcybA+LBhDskyoJQlgZyi5a9cbgD5FM1pF7quIGB1TYvFE2nKUgM
FsEmSPCpgy01MbC4Y1E/NLsFrKvfBSDSeYHp5T+j5VygzbGwLsegwRQf7HlkzbbbMhSBqpSYVS8T
HTqZKmAp4SI+T1HI1a/QwgfUNfxrPvpqLhYlRaUjPW3HfiYhth+TqsvxytMy+ZSBENE52QjTP9Uz
yoZRxDBlMKwTGWgECgS6KgbwH1anMO8aGUEkeQr8M7qEgHY0eGVhY9kzc1wBKLiDLZyBBy5+ca2g
mQbVfemsIkd8a/byuaCKq68XuFkEseZuQN1os82NXWjE1IJN/2n6esn3kGZZEh748aGKfNMhDvPP
coCihB6yBB9ZxMSFieocBa0IWFQwGiRVk2CFpUYsweysaQnKJRcTTJr+1cY+5o8hkmGpVumpBgmE
A73guZxIq8CJJ7/Kr6l2jdO8Rq3us3KKYY0B+onKKVwADrtYMJEsIe/SCMMxjR/0HlMaAhZW+xeP
hLBb8Xo0aZQ/HrZapZhx511KmtY+oFE/bZpD8Ns7nYnm7N2VDkrM0gtldYw9UVm7hD6Z49vyyFJD
A2PK5uCf2aX2MVt0QqZYnZ/acR2lrwqKDUgdE11QEx3l8RAl6rPu/ztLZd+6xq8+GTfjgb2WvqGZ
XCW9qdKgVzTAwsLJqQySvDgWc2vKbmyNrKL9rU9AQ2GrXU2U2qvX6pTQmrphkacUERAEQg8/EO66
tu8fO1KegNHsObvcNRJN+nsUbb1d8M1Rt/enFMmahvMYV3IW56CERSwR/cvwR548+3HFd2gEeHdR
3oYeHOp1Nkd6xYtyuJ2sVbjnQHC69SYEGwt4AW6l7ppOliwhKfEGmU/nPMXrPtMw8JTEwCd/o7Gz
rOgrLZtEBHipyETCSfQidH9TAkhipF9ZgHwcq8uygCHxNfhywMsS7dQovKGS+4E4QGGLZAzHU+UP
q5I9zT/lDYOobF/mEOc6+dnLmaksnNp/EWLshxKEupAh6CWforeXFRFT8xS+J+n2tJ8olhodYtvz
Wo2MYMHKVPX1c9k9uOqfaCGQBeRLqbNIIL/CG5F3B+w3EMsQIoGyLhY2TJhnbZqbrNMWvKw7Dh+G
5nXvcRzkgyvbh+bo7Od/4c0e3Eh4Rco7Zvbb6pIw1fIEAFAUJBmTZS4MHLZSgADsUkRpfc84t+pM
WbPWdRZ3RMCLvxK1HeBxR9ExV7aGZFdjkDcft5PmtfxvW48zKSasfrgIf5Ec0dA2EMZbNMuXwPdl
tgM61zIyu2FmSfVT9eJZLrc7KgHnQV9gg1GONgKvHJm6sn7oyZNs/EgZq0c1A1iddQDU9sXI7dWm
HmrkECz9bfXqRuD0FHOamslAISYdA3X2XdIQ9RStjGZPOV1W1Pm8oCnHF9ul4aXhdgTaeRrYuZTE
cmy6uwnA0y9yspcKl3P0AbEpNqqrbxpTvEMmcCFE+bRKFfw1LGDrxKwAbd5F0CswYvhR3qnnmuww
AnoJujMyl4upn+i5EGjr+2z0HjfiNWgwpZGVxM/+sUmDUkvT+iVDYGie6pn8XG5IxueBHbqwwEum
85eqeuS9Pz1hBt8ZVquAO1y3e37DB+FRlKyjHxa8YzFnmMUeZDacc/wqK9OgqN8RsYVqsbw9kyMh
pP+qCLnP45kJ15+pM0eDdoIR5Z0vasXwO9gHyX/K49gwOy/Yj47A4HkeEJgcWPPtWss7SknJHkjN
rcm3q2fFbdhPXYfFj38z56ijDUlfyiInbjbtZv0OSvOIuv5ftB30ee31TevQH/+4tfCV0Qafu7Q7
EcQkCGIOTvzrpyCNVBUxhGm/UD6gnyE2cbS+ibZc0ATKg7DEJFzlsLSIwFHMhrn6ADn4BIpOs41z
W7Vf9HGd/xKfzN8w1Y4TmfXuZMZT1wz0vMd+EjnII4EdrC+mNXva6OO3zyEwFvL0bCPd1/3iAxMz
MvqeJ881myVeEzZ2ySi0vQpYfCM50Nca/KvbRLzHlgdgJjUaJ5jj8JF1O9v/i9OvWGLFS0ImGQaw
UNXCs67/L3iAdu+jH9XUTLt4UeOUakd0kGxpXVJdGkAFgi+ItX3TLyRfMUpdpxV4g1Sf60yspkj1
bdwu8LeZd9O/iy6fR16lFqk/jde4NC9njdmpfnWs6ERCWGCA3z7/JfIPuOutl5E7RBVNlNPvc3d5
uShZXaN8Ek8p6Zxq0r5EJasW6zFdRQXqAmiGlIw0BNvEFPenCgxwgpXj26qg+JmlP81Y524qpyyI
b6ezeBOPIhs0xkWuwjBG7lT74bMFlVP1f7PzCfiOj9PGOEmE7n3feUwCx8iL0j1cLLekSAXqbUf/
yeAOs+trSsiKMPAre6TakdQTm7YLHQA8I4LmbhTDttfqPgIT9aZuKe745++D5+Z+iQbidi9OrHzT
wlvlf7hAWQWvWmcI6PYuNiN3nrI3qpslzfqVUEKkZ4bUaoCWGS9lajM8RlB6BVn2nl7X7HscbpgV
8O2NwQmn04+8qX3leEhB2N5V44/mWaJi4N1Sy8HHCAQuVPgdK7o5Q9wXajwg6Bg1aduBcydSsg7N
W2Z72XC2XSIYkRakOk0+k89/5dFyqPMi//Yr2QVNJ2pFbN9pi05iDtDyQwlMP3KNeQWIk4nxmWPD
F33qPicXTvwUDpJWsl+CyuMKo/RcXu8p1PCHRWKhnw0+kpZqvgfo7wf0EywiFYrmSBJ6eSgfAK4R
SMhjiNqLFXSTSIP9p671yCbfftR9lEzWz6P19VFhKGUPx5cO2p0Eeqj13T6u5E2JRzwjvEK9essx
1PS3oaXzB7O8K5oaseF94knvGPG3aESHbD+xj8SoH1xVPlzkeAXOlzI2a0+5X45KMrCOzrVHlztH
Q2d+Hj2PsI9sQRxAkgg3yqIoGFLjTGOqRoiUK6YNo5HUP/7I0yP47Aex2IWubNwQi1vtSOmUh46o
lhBVhrOfWhHO8umIXmGx9z9ldHLZTA6sgNIKU61w4t+0uTje62cXnPrZFvAWLmosy8uJnfkQDb4u
Snnk6atCK54NU97adXP0qiyYo5l1fnwWCzV3tR0DFchEyKYLWjZmECPRcW2KoYIPNkA8z+Bhf4X4
//ARC33xDhnsswqQPAsyyMgy0SnrzTDXW/MWanQwUUUey0ige/mGoM1iIb5tt31U8aK0G+3UIN49
ByLn47z3VmtMY/lvSiMd2pY4enUSCXYXvDMFrlg27s8eO+QvNq4MJYh0+RHQKCI/xTswWiRjUWkN
sjL0R927pkPvyvBuZ0vCfs0uvCF6wlSxpc9RXVaFgp37l1pWJdBoLi/yoZozvwl2p3XKtmVLG1f/
Bi1jmoVbqrJGBZl+d9sIXwbM8fYca2no/Uj5MQIi6+jcuq6DcnJKDT30cVLoZ/JQYA+me8uVkSXQ
ZKIrfErzANSebQNzEPux84oAFAg9RkA2XUmRSV8IeF9BcW1Ls9YEOEbXFUxJZauZZo6FkvrTRekw
Y0YDTCwobO13aGDRMDSQm4LSCpm6yfKLXB1qm9WcdTzH4WKuXWKgiik6PCFEkWqvu6XnlNXOzz8J
EbKrLZWVzheivLQ4H5wlqT4WEI9CRh8Igiw8kypSP59m1H7okZf62FhuOormNLlGzLurfpPs4Y9K
VlS1CIxW+3g0JVnhjJTNaUBJLS9P/SwKdeYFmL3ICUURD5/6Q4PFNGJa6eQvyeFvD4hXBQXBdTI2
DY4sVlHOx8LnKCQZHeWqrnVcdjo3G7YzjF+aOEJcpvjMp3Ys3RgAsGlDGqRQWmiK3TU3HI2Hb/e8
4RnPfVH3MHKHkAE8Cu8Hc/S23jL3mPQNgykeFIenLCaom9GvAYkUBugtfNSCk5+2WJjgU7rXPjMY
+G5DtEXJUUaVYuqhHihtaB+hh+pAN9D9uL98DNz5kfY72w/0hZqGWGru4uJ+H7z8VjBQwY5A0env
NZkJLEs/NT7iTfsLSDuFOWKNOVpUlrpgIYMk71c9hs+1j58mn0/5gknM7ZT3tXbJou4UJtGnT+lJ
1S0zDZuZurLhutmNaPgP/PkLO9XrFYP4Hx+sNW/3EpY2LjG/L+QouTJ3JB5vxbjC4D6Wn6RpSV/e
VqOtUZoeiXG0tBoJGySOYHlGcvmCyggu+ntuHc+qY2CxmnDYxH0XdpIAQprSOc0w4+nkcJYwS9te
iRDR0Hs+Ycf4SreoNkEuSbX/MOh4S82d2hsay/1XtkdraUKl4fNgI7JVP88zhPJOghcIy/4Lq0K1
oCTJI4qRIRh9duBmiCTCd8ghOHTxneok2dUK2X31+mdpHO+3//8vilQJmwnWItds72A1wgafAIF5
qLVFm0/aRHEINRLKMHaPm3Zgumxb4nBQweUWiIfWNqOOCQ0zIZMcxHlyH5EE97jWp7BKq98FwSpK
ipQpUys+5gwmAeuy5iv9kfJCsXM+7HrE+XVyP0auHDsNetw89QDNDOXW6eVFJFTAN+R1O+tHNbKS
qOeXoGYfNTCQgOlQHkRpUYEWal/r6lX+NfDANeo/ZJr3JGXiCK3u+5tmxzeL5RdejSFvQaGBnVM2
oDbY+tIAcUgn9JiRFzwgrPZLvypfCWbtWWj3E2NVofjLgKZs5uAXD91f6o0yMvGeUH8xY7x0VyqA
AOrv1nB3z9TyAgmcynzJjIlJggit1VaB5ke0Z63Ms6Mp/w+llVHKjlAB8OsDNdLMxcylv4fIZr0O
SKqmTcRYOEu7/KpnyShIyZkFqgRaRbtjBcz1QvWlY/o9NEmAgaluSziQ0UND72Q91q2taZjXXjYn
57QFE/pdfrPFE7S5mgJvl/iyB5F0vZVflfSu51otr3TpcC3hhgp7UqFLp0tPoqbfjp5VFdY2V91R
MFwdEmPqzXATy/Y2Nx7aeyvdoUe7IvCzxkTDs1gbvufZcHA3unJHJhzE+UFIIxlrx6pzE8rYm51s
r2v7PQZXprp7PKZanmQODD6V5oc/GHPEejJOZF82fvX1LlDDWWUPCuy79E05YfaLBt5Wag7HmY6Y
86vhy1gBYnaWF3NeGtuBSmpz4qtvLu9/uL9FoZrbTh18iwZkLiCGz9b8HLicnDNjtMbEUm2SX3QT
nEtdW/3OBB/+PFL/FSaRWcyblwQV+mfpkdJ+dPJy+wxu5XIH2uPz9H/qtqHVGaF36U5YTpr5c1pG
4u0b7UoiF5yX1mVRVTdw8pPQLznCsiNpvKf+8m6yxn1dmp7MuScgeCjVI5z+znHbQnOPK0Oa/VYw
ay2mIMpQoLfivg3LmG5+BRKq4nEsy7SIruiZqTK8uThUU6MPcaSRCkOsEjzjpAo4w9SN2WjlVy3g
Fm91T+tfh+2QdZtN1U4xBV7KSfadD/DK7gOX3zfGAxhkQfsG3H2xZinC2AcizVdanR8334eYxnV9
19VcA49oBBnh3LXhJMefe0SE0WDDyYRezAK6MZ0gka0mh1Z1oCC3dX7qZcRpFZb8G645X2X98MUS
SAiu4REj+TjM1OokvZAYh5LKOL2S8nSVmZIjodO76swMf4PCKq3ecs/Eu3E7sKn1WaYDQPoeHRAg
e7srQwSKcZ2PjDxzSOlaS7mNxAzwPdHca1OhuFaFZqVLf1spe8zYEXBlJDPS6tH51C70AXbKbJTB
eDnptSqFCUvr7Cw+1S2EvmgKsBIrA7dZ4juz9oZn05Riwsi09pEjoXQBops8+bSzyu53id4xNqrC
IMlpUKmqglzEz1dqTR1QUpFpH48vvisCwPwo4mCLYhjabLP/u9hKQtGdtiX/Dmwmf/CvHjELjOYP
ob2YyLVCGZTxKNdd8ccWJBcXXfs4NO8qPf7/tFPOVtOzTCTthGhm7a13Im0RTQFxlYlpLZKi32Mz
Lh4lzcC/9BkUx6Lwv607QlmiRVfT9xixLqUM0DcllP/K8JPCRJQ+Sk09KSMkUszHYmu4qEjmfuLS
fesPTDcSL3ioJVSkSvrRuWao2oR0pw/mBLw0cACOym/V9shBdQK88MatxMvkUEAf1bCFx3yCI1Ta
9ugWcmznR3y1DZHa3LMBUrAUuJqUkgs2dltO81aiF7i6IigAshrauhdwbFiYsWwWUOk5W57hlbDT
NVZqricVxOw+MQ321Vd3B2A8qfz0mrPHjG5JYXDfhq46vFlyM0/xJ+AOGjosMoLcXZWlFmiIT1Ry
9hh/IaEl0G8SaBF4tB3S3QuyEDtdGX/pPo1/YgF8jjoifmvBtX/A9BOfjFoFP3Gvl88M1TcmPpJN
+nDxJi08ozeJYtu0OJEbTcp26fYXvWG5gS5K7+hGs2givXzoCbxfQepYeMBanaJz/IfJoHSYOArk
1ALNzteTC9aAVp5pPbHxfmJegsm1/PZ2CDDvd7aIUKHrQcnnX8GNN70mG/Wrws7EPak3e7vNqrqC
XM2osg0RBD60h47QaTjprz1SM+9LN1ejVQH2/XRQWQxTJk67Ln0T/XUNtYWqA0fCbN12mrUY/33k
nAq0wt0EczLwSzg7PB9d5ogbO6PG9NRCu39ZCcBNKb/A9omawrjopDOA3IP1Sa3em5yj6Wnq1euQ
Kim1Iyway228xp/AiNxBr/iorBx4l/8+YCMp5GuO2oYGiZ984ClVybJ1ioARmKRSIjR1AIkQYBsa
babGwmDGH9etFd2m4/sLNhKrHK/PTCmgSw+Ewt/vUB/FUxYg8Vu1vw2SyEOKQOgl5CmjJixLSvv0
Qn5YsK4NeSogDD5b5C9qE0AqrfweiSWzAOlEFuwmpXOcRmEdekV6QsU7N2qTvFEWZ6wPYSMl8FYD
5fIMoSVVKSF7qapZdPV8+UuvqAfsAv5kw19zRyBS/Ge3kyA1hcQtXWzHBqosuj8Z32CFgk7d9qnA
Lhz6hacJv4PS2izoFDSPygKDhEAse1YhEPVfrwqLcd8Nwa+YNFulWpuLTKV6kLKdq+1MCKvZhcqI
AK5RIzKzEiToDCoMGm8HhS8pqr7NJU7Wp/OGF40oSgBToDTG/XB/xgGcfdH15UwbDg8BRbjJknHY
lejCnMh6aUgB+Wi6jv+CIQjvF/DMD1S1Wf5X6GaOU/k6iY8Le97ONR9mlsZfuo3gMLOdcgSi0ENn
06eClt29S3geLCondftUg3voP2jPfuLJLsvMtUsneft6mC/9WKim83P5XWkQUPiSGa28KFewDDl8
KVgQi0zVDS/t43u6/eN7u3z9WSEP9NV/KWm8hPYF8zeyg4Dvm24pXEdOg9wb51lecSmYFjv5odHP
OlA3MHPvlFC2Nf7Rf+n4YjQVt5oR65YPtAi0fJNpEEVffQhNk3PsLRMkEsBNYnowUV0Kki+1bi/V
ZxTHp+LIxi9mU63V0Ivp4eLO54xZ3acxPeOP93VQ8gAfNkng1JDOSr/JGnwY85WGHzSSIO5MFwJl
cf5PnEfCgov0X2OgPAV22EYWNCv4BdF803DMjFj14/NZYEqUstK2ZEjmYmNuPi4hQDVg5mjRgnBk
HdGp08DQ3Gl44WrBtG/t9b5f5JjvZbzCtxRBTNh71QSx9fbECIRfLpU8HpHtcNlPJ8igirrDHrXk
Xf7lLEUtmX0QYQTx0fSuViriXMeOKvg5J/mBAqepfv5C0ADyIrNkEp1sY8hC/X3wqz0m4RdQDZIQ
yOgAGrozLtbjOpSwjrFqLuD02VJNFoqWnhYrY83vQGizrZq04KVfpdkJ0R0R6dFDWB0I+22s0Igs
+21RHDPEHBnhT78R5Y2DnmM3RBEIXuyjq+XLLZJBM6wmUuRQcjNtdWGPd6DzajatfFJAH3hlEToI
ugL8PM8jWONP7SBi9RxAzs8RfV5FjvmktGdSwSRaabnB6NHEl38RSKlkDFGjJvjeAs6cqPNS9Y6u
LgSow8RtkkuIkeXwey4gvHw1oHpQq8//rEeaKKg7E89A+tlWIJ90/9AGrYFhtwpHIGRZm1P7621e
gERW1tUNDhBg6V+DX5lurQbxktr3gc0CFTejz8DaggPkJyhLSNjtKQA5lWL/gnzWbcakYiN1FRk8
rzhyvdgPFbZzS/97zClJiezfWpJxuJR1IZyRaOFgBBMSPRERnl5kb3+YCQRE85Tryh3XGO+4jQgW
UOcjKv0jFCBr/HGiIK/pBEyTJo8NBwuRA9W08vTseoJM9swTifCnZIAQn1vfIdJEVlIfHi4rcqB6
OqSYF/ik4GMJ6t4yv7G82IK0fu+TcR9h+0OQMLzMKZR1uPKLEk7XBnrLOjSHRFPpn+qENiDbYTst
nPIkquFX3iiU0LYRdMzceQgw6/eWmvRURS3Vxnmw19MbQEqJFq7T613b45ZwGky6YCP4er3LNXA4
vyKfRlIbPD1K6ZTmq79pteymcQKjskkYdZtXC2tQWA931XGYDMUZBWCrblr8UHBTG2xpN1jhzDFy
DfU27HCJnXqZXyppnloYQFFbYBIiqCcALxaPZiHj4UtSuql8mQq4TEqNpqnLhzA1GnyiXLep5ywA
/gp5uxMMbZCedfZCaxmPve2eazcZb3QoFsLP/ZDnIbCCOvtXCvrb9Bu/RDjyLTQBxyjWihU4hpsJ
vg7HjizuxINB2rjFUkt+heoga56LpkUXfgOMwZDz9rFa+bzeBgwAKT0/2MkVv9VhkgtCvPIN19Tn
pcPlO2MwsPIqvJ1nEvjaOGF31zYJnp4dG2i4HmH7+9PMtg9Jd4wHZDB97YQTyayAyesK+odPW5gj
SlQevi1oZEtFcWzbVKfMqqV61TgGrDZ9RGB5m1JSMDIWgYej/9a4G1gHyVHIB4brmBMxv+6uR67x
35aOM4B8sKFmgDZgLTLcVdP+S6DG9tvFWDNYdc+Bhex4DW0nvBAD+Z9gL8OaJn3KAa8OiyMc1Xm3
ww7ewxhB1qvt52xiCYIiJs7wpOmL87cO697/LcVuFwiTRYqRrYQsVLXB1cgIISH7vtHNdVAXart3
cEQZlxd2qMTpqbSX00pXbFC8++YngDLbjRYXBYroSCzn0N3g+ZqKNiJ8h5l8V2qJESp5fGGYMR/p
DNoxZwwb+iD7dVP9iCB0SRfVaqJ7w1TXAfDWpY+qAwXw6CNuI4S8XH+O2/h93Su/1aNqc6+X8rR1
G5YYiPgFtLeBpmpVHojS+0U866tde3J8bmZbe80kiciAV3BzZwO7rppGp/tcO2tJahbdwyQnk8Zr
ELisiIj/RYvDU71E7uYzPQUma9K2PhVCuLp13R4MFCt0UtSiWScj4grsXdEkKIWl7BYC2uo1Xot6
nzl7eGcwu6vjnkupBHKnT34DvkdeDanqXSPuQfxGTMp6FP3aeQgyySzFRQTNWbMLWMfvSUyObueS
/dqdi9kjKpYXT5hulJNeyCZcFCt3wJzoZzfBaf7OLltjEGVuTe4R8ia01jW9K3pFKAug5yy906x2
vDaroPhtFul/XO5zs0mM4qVdAeodU2/Va8hct2leIcxKxer0qYGWua2/JJwyuap5ki6L7TIwv0uG
4lAVoJ57KZKfPD4ECKduGSxRHI+4OmPkqHgdMfsm1HPOc1TNsy2LbK1pnuxYYbFlvGXmc7aUta+W
w94YIBzciYd8iEIB4GGeRf49lua5MQZrMmbb7v5Q4Gcl0TjgX28xaO3nz4wcydtci4/gyrXtWYnX
GbDN3IacGHKRjXpsgEQh5hr7oIgEXcDrMfz7G3IRjOoexEeNfuzGVWcMSt8+sC+BerSyG4DIx2oQ
mLKo7ivb5hkrfrO+oqgQPgKBH+4H0n0HlSp4jWVMmsfMHeZ2+sAq5541AZPgDa1xNcsqrhlDXcoF
+3r9rXD87XL3auZ1pTw2q31DY3TNFGgoE3RGSrchH+yjRK56KD4NT9hpOpMod6PcoBg4iatiqijl
uLx8YPp7NU0a45P28UDkxABKmkyO5dJFzYxNnqsXu9VFj2R05yjQCYdiihJWCvdHNHzobWbqjOZg
F8zfGLncVktNq+SWvjlW1AQtsOARbCW6STNhfeZ3F4kh81+Zt3onbgExcAY42s2jVkTXncTpNB8K
Sh8u+LNryd+eoinA0ZclTVCkKcV95N699DtXV2MkIeiNcLxOq1Se8OUyeRcMyFyHEqeh5yF2z95Y
aC8uEt45RFHv9JQFMQn7+10IrE0cpekAgEt4muxl3N314jyWfEbSfXhfkfjIqnYgmHldog8YqjP1
hBltdY7HcVC83+RKPOUzW9fNClMSYV9nAcodgGWIZ1xMmrxBrVuZi89y1o71iire+Z63GZMgeWzq
1rkzWxVXkVwWPxEjVmSTa6aonvLFVy7HsDkqOhWkixqT+52ExU1doVbzWf4UbSIsHT6+Qa+G3uat
8LVGmIj0DKaEHaIGTs8cP8u+z8PWqZUZyZuh0qjd1RD3Lx7qSv6E0znPSNJMyvnTz+6w2/OMohtq
GEm7KTUq5sh3FFcr7Df/TxiLY6ZOC53NXw6p3iNp4m/+Xm8yBLXdCMDenjvJubgthjq92YMEM6gx
OQdddCcftHkc5VtmQWpFw7mKRCPGLPn7iKOgahPFQL2Cl6XIi4jNIfuv+OBNRzlDLhyIW6RtH3Jy
PT2el6XLjr3Xax2cDL1npu+U7PzbWmC65yJsohQ9Dh6NRAYuvzgj196R1QERfLspNStTfzBeIp2E
ybmdJXaO5rSi/Imhx26xmznfNMXsDwr9KhOMQOAdtBnDDw59EwAofIl4/udBrDV/fwV1K/l+GlFp
Hqer2vhZZS6QGO9V/fzduMOUaXXwhOL1ylG/CygC5WVIxJtlRIkY+8W3e5t1tlZblpXAYJAXRWIb
gDZ6hrzPIG2rQrlVe2f9w3SIHaOGoeCGtwo7Y4jJVbs1mdzDxpJUI85nK1057E3gTzTUS0Fheylm
C1wyDNUNFtGhfO+cDjDtiAUzJxen0HkjiZYCR8d093bEnhMVGLct6bdw9NHcmjd5abeH0HvTjA4i
sAue8gF/YinuXqnaosV0kbv9OfwsvUreF9Q+V7LCPImj3jspwiDRP9xH9nfBpRsIUpOV5Ixd9H2o
nzAVTZKDKvJokpJZXPQvjU8Ow8GbCUvsLOladUZkakPBVhTNQsWLgSfLs6lvJ0rHUCYoD/1fEncQ
5JsA758SGF2tF2U+dzLoZMTml8fQJ6VTUvKdezuWhVXZ8KYRZ+7/9Kl+DaPB9Urbi0I2yi1jYDbw
krU7QE1BNgknZIaDwRhRbBCvk0nj9BaGFZsOhtqJ/B/IlLcYIjE+yiaSrGu43yuTlUg6ZTWYKhoO
2Wd8jOmGLJourO2Pwuo7b3VbWchzcuQAOV3fRCNulMFoOzfQgT6mo/61gtGHXndKuu3DTvzOqOpz
2bg+1T51b1GvwAYnYYVa4H8JcyGUM90IOiIb+3tsHZiL+zWALr2bN5RW/p/8L3bVWdH5fxfWxJdL
4wm42rzBw75dvkd08snmXPZMo+hXwuT9cFFO1z1QdCJWShC/pCDAIK8tmjB+gck8+XWfxhGTz0t0
kJI4xcbhYL9+/umzUz7SC8f1L7roGJ1Dm4eK4ngDd4qewT00O3fbXDMfbkL34Mb8edcUBQTE5OGk
EUsHelnKgkmW6/259S5UZiMHoAWnFl+Z081F0xFaq0i3SwPxQE8P91EvpHVDJnexxt02Q4/Hi10o
kYovrzK6JOHGII2IRsJy/JzlAqYhRVXZ3Z6m9zDsyvCMA1xEabTyn+4k/bCVwfcYOgJ5W4YU5VNo
9b5YdeEYf72sbldm1gQ+h7nZhLdYlYi7g8aJIolm2LB/01PeaPmrvG8k0iR3T5xkjvQJt0FfvPSQ
A4tb9VCzZTHqYNP0AZ2NboZNBlR0/ZKwJ4ZNl6HMmo+mFzkWC0u+C9Yj6IsL+rWK6ql4Yz8SD8/E
1qzGUeMP0V7EB2Ro96gQtpURgnOczD3oLEtnEVUfCBzzhbXBAbAusI5R11jEs0MrqMME1WjG1xFC
1EkgqKN841MmmHwivmejakA/LLEsgftwlEXQSGyu6vsb194KmMNIXQzS1CoM0GySb39OedxBNd+7
CisJIoY4pInenCe0nqmYYTZOjd+XsXYYmx1n3VMizXdGonrgcKm1jN+G/w3KBEGFmsxmWBISaqgQ
YDTkrNkLMBPBvdknptRD0OVU/7BQmaNQb8oVtUIRFk+EWgz09iWrWngMS0bF940CFfm0usMtKGAK
T4NIeg+HOr76CX7oLD0HxZK4dsEeOLsDOBJw1yZ49rA6QjhjvHMGfoJ+GsM0w0tnEspamX2ocI63
g79U+NtZ3JJXSrM09C3fq04BpS0PUZ9DoJg7OxY0aMjjlRJ9rYp1r/8L3w5gvnfzEcsxS1qM389S
8GcZ7s1Q431Bi8jFpKFBeADacCvi7ndwkXqE6x5EdN3M7uPPdxl4pY/4AKrV7UVr3esnxVzANl7E
P0PW7wDiID6fOls7cwzteId/HrQGnkp/4bD+geCMr4/BavS7SR2ZeSUKhsFFSXVBXATtpL2JUx+5
ELsGTEOSUB+dR713/lYgElXSElgKN8nL8D7MlHY9rNyWpC0ApN8DiAxYO42NZXZLSNAyOO3OpnYP
b/iUEDx4Eifp7+F0ApjJMV4mQT0gjQ/1ZmLQ8MdfYmBrmQAxupW6Hw/H2FPdg7kFEdcVRfTTlsc1
rikfAbEX4PN4x2aIVzNAD5fz1wHmpsBrooFOtd+714Q6YbWDSru3yrYGgU/j4q8apPS7dMd7PeVn
fg+i6+/sWmOsKjA6KU5aw88qBKuapTL0F6vDUcT/0NYiC32G1R26QwmJGCZ++toUFmPVe5VnUdwr
ZIvC6ky5Sqkg9X/HrDzgOX8CJegFqzo0mCDi4EtnRAK9VD/t+3igYngAl6bot2pgyXH2cb41BaDw
NGCaSu4BviwN6oHI20hG/WKbl21KetVMhagnTfX68P6jqNkHOvR4XzP1lrEbYmw/GCIjjVVWjUGj
WgzX3gS64zIRtS3QVzLsU/Sxt1rUWVpetaDIYcVcLFrv2P7bxbS4IfsuleFQxjq7m+YnRZiPsRrP
aLaKy4QmnJxn4EC/To/0RkDG6azr47ex/KPg4s5KSi8am6fHmJaNr2KDqngDYa/2uWO+OSmu1TAb
4wnL1K/wZdltAa26zCaDSnBpqJN4rQXhU92tnLpgcqT0qGtCOmb2n35eFg6eHjaTRqtPX1Ucmwu/
hYbHI7akFJwBnwrAo24FK18bCdhYk6OfLtx4wfn6+/+Ib1gL4qFbSZI7FhSVLSNd5+jNfcCaGRYK
YymvNB2FRnoPTKvN5bgQJpAznE45BcNbTmvfjkaiGoNg+8mS9G4/CRg6IdDNQHW8PylgbWUKhiM5
aMb8U3TzI9jYgX9iKKME8nyswdW3YPhrwqo/Hl3TB9aiF4/wpZt8LzAJcUCfttgtQ9BHpZMhvz0H
710vixp4hD57Gaqwmp0+BOVDE2128QPp80R5khoQomb7SBmq4WjDjdul8HVk0u06sgyCpdPhy6nl
lTcl4rw+eYRFzQx+TlATGxe7EBMplaR7n1RHnmH7S/Rpp4n1TSmrjfLsmCR+kE+9GmVykL0XvT/i
sgE/D2ILLi68IfR6v3/UyoAsIhZp5Z3D87mec1ZBsWrwI3+m1jNCv6sDGkSJtH8acYzTZxC9JZPJ
LQgfZnHQ+88A6KjpcnSNx2D4TAAu073giY229qlm9MczISullpmRu2OSOqC5Wn4Gy0AhpIwFJIeA
DnGN1xpKIUHG4bESq6okurpMmNMvTLy5oQj6+lFR9PHL8qjOThAo5w2qOp1IECiEFjQf/dPRp/vm
oAoDy3R/3CGBjtIKmiQaYaaUGp8P7QNVyI+zGw5ZALcmeVLv8tgrraQdNfS91ryAmcX5JQXed0X8
gXmATiO9o1WCKwuAEmkZh8GLIqOCfbW0xt7BkJ5kYtTVmLN60KuS97oMysbmXQ6LtZ6MPhgJZaAd
fN7GlhqWwBBNZeqeNDEtyRa1xCGsX0OevCR2RJJlII1PnSivk3o17jnlfD3rhRDlDtrUeFbgyii7
KoFHNHnuVb44pa4lzcLxTeBzby/7ISx7JiNh98lRrMF7A+d5cpDP0ZTBHzydU3t3S7sRnP+QlfXN
EqgIepJzZqiZzBHAiDJZnkj9/ZRHK3eJORbo3nr8NRz1iDzZZRdVYcbR2VgMvFH9ttwcboZTXAl7
DS/hj3hEMHoqv/lPQg5/k0Cwp+uMmYhKIZxgMUNtSDgKexcGJjyZaA5XVde4kCpMR8oX2s6oH2zp
Xx6XYVbiMhcI4R92qQinouBraHYsVkLxsl64TCUAmkIuJ4fqEVtPvWKaAJjT6j5k1DQFNtlcq01P
h61QoeyIHq1Xb+B+lhzvF7jlYBZpN0rr3dqqNb1DATlPNWsqZ5gilBfsmVVAwQ/2b1/Teex+EIdz
+1cZm+WTQcmkRkO8/THL2qTfAy+aJZrVwXIMVDX0Grz0wJe2+FCYPsoOBntitVM8vkHNOJH+PsJv
ugS+BFl8dBKrOxWr5y52blnVefFO3NDdp5Uhr7m5ON/wc6tkaPRIoF1qqhzxEsNJWP56BzTab3Mm
fwMWnFlRvcT1cjGqMH5BUF0ZKGyUeuZ8T0yxGYdugB42WUAmCVWx8NgdpF12ILDCQUqgyoG8tL16
uYCCmUTjwhNTfhCnEH5FS5auHjFETAg/HJJJ1W5JRWhvYJZe6sBoeSBTi0FJxeSne7/ls5syDZlv
XPinqBzzoNKPtNFeH063IPn0AmX3FAthzkVIw0jHh5PXXs0zv37XcEYEdR1ckcwZ49iyqMIWGHnq
CO7QJqG0wx2K7JU+8mWuIEWCENl2NO0iaqsdyKqYpZx1g5dYvt2AnrI5mqXLm4aMr2uJ7pDELS8z
pnb8+j7J86yu6u+lZMH2J4m6i1YK6zSjrYOw9oKR1ydkD9WWhWoXLmoooHa7ziL2gowOBY5iOBq/
0gw4xIBUCVSgXS6cfBTDyzqJmbvgl16iw9tsgTrc8yIU3zKNGqVbeSwRhfZ62Qs3iZuE3l1Pt2+d
iacz1pScc/9gpmEWTY/eY3B5+TCG0ku5e44+D84O++VLQjM970qitd3ivvRjO65pUuKd5L9EkeQy
lcC0pxDy6yMHJvloi2HtJpAYgAfkn5rbtF2feZFRYW2y/ODSX9hSdYT5jfCqmyjBaEBGiZYYymkN
nWZbYodgddfJ/duzJ5Fgn/uCWCDvobjtb80UX/qkGQSWNGhJ2LxRG0x8yAK8u14wRXOHvzwxs2qW
LDJslMpDCp+kxAimglLXCupPzdJMuO+63SYOMsm1plSXrfbGvTrMS+ma9GsLSOWVPkwm1bbM4UzS
UMHwnbHpkl6EM0N5MQfR0HO0E13tXtqKVeg6HBCO/r811Aq6SCSqco7zPSPbfoM0T+P1fN67c47X
uWRTNRSf3Mh40RFnYM1roHdNIEypRZ4RmasekoHdTAA4JTGMrD1At1XEdJSbDs4GhguFNsl8dSZh
N2n14iR0gB1moyvFxLPi+3OclDdr33kL5s6lzielas2XSFONsuw3mzL6VfgGe+Ayw0xlSIR9nQGM
bUr78y/xXAv5Y8xRu2nU8ZFEs/pzlat1gelVYdUrdT4m1lH7M4SBSv2azGLSjZsX0FWO+leXBoKn
RiR4wV7rb/Vxip4FwqL4alpbDgHQkQqf9hpUJinnYe75GWlCQRGSoYDU7TshB1r3oEpXB0/CY/qN
Os+4piP1SImuFLoINDT3dIZJs50yeWLOFKP7b4fggetMiVJhbYLzn5L17nvOczsZ93TJ701Jdx3m
wwEvJKcwkjZQXsWPx9yuGQpMsC/FTDRk2YTy5PYdKEwx9qVakxINVABWqpTS7OoNW2Ei3G5Eu9sl
QmzpNona098fKeBNghZOs0c0BSbDXSc48vyPkPGQQ589kC0vHPvRD0AKH9NOv9IKlSM9mcFyMV42
t88RFAyMb1nYnZLnxkdtJgWXhbOxgUg1ywT1yi0Ik+EBUSaGhOnQbal8M1OYSY9RL+xDwysyhaRJ
ujRbf29m+xr5PAkhH0X0QOXbeHq18uEq87N1/C14GCJb6lLF2F0OtFRlgOvUkMdD49eJv/J4WaN2
sCOdmLe4EQd6xQQHmfSnX2tYXHEYBXuxADT974hIHPzK6wxnasCz8050NYhoy2c0MEjlNMK+3vO0
Q+0Wm0AubAabnJaemXJEGk8SWW9fDLjHsAojknMBtXrPoMvnQ28eg3Q0aOiVfdJWwfGM/d/od2hJ
7f3hr577Z4a2eu7ds3TlLFxX0a9xHflCQesIF1jgdKpaWVulW7u5LK70J9LA2RBbvUwwTHSSKVYG
vd3HCS0WZHj+fpwgOggXSCZ8x5L1JwcYrVKQKXDrWx9oCNV4I/SSEqgzm40CeGckJlbO9l8D3vyh
ZkJFK0eoIEcmu9ofV0pTFM/hviOC/t3hHqioTgeSi9YGqmPj/+HSMTwznKqkMP7S/IiYYLVDA8+6
LgM1oXZ0rMOV9Grk6QFz6ZfgJOkr8S8MprslMWpaCPpyhjQbeOFML3VRUdz/sewzoLtZsG5OWmrG
6hcVk4K0CvG4voCKEUabjAXWwrDYtiSZnVz9uQfNpxCjvQqIelBDZCQL8QFcVgxLSXutYNTihCo+
h/pwBMyGQsAU1AgCrxHj/oEA6eoIQ8vZ3G1rXtxCxm6OR9eotBoLzECdVB6WUk3pC01/FDs03xi7
+yaHD+ZjrhtPLMoStlsSIKlCyrKISwxoIwlzEQRngaDyrIlTV8FKvDX4Y2XwUGgcrndgqjPZfeGZ
LiUYZONYn8ELLy639sm7U2z7WebdcGkRmiSSN4zrCIV6FIKolvQYWmw1jcxROqfGf+2zQaRkf/yp
zd9i9XMDCyk4FkYaDz5FP1O7F7rdankFeefv3u1sEshmrXA0tOQv63weY5d08cmuHIk0LX2bpt02
KxFgj3cuiSiLW0qayTHqkqY7nOBMYmh0ydS5BzQMoLGfFr+T6gPl3duBfOl8UQBV1UMg3vQMwi9c
KE1MXJ1vyVMPS+j9MN/8AISZ/b3zRwRezq7Rh2PXJf30fH3q/nMHE6D5/8citY/Ysw+HmWXGtQpG
IZzQGHAmFr0R0IH+OOWrgPAW0SD+1L4AhcAspsBwGByWCoC9T82d2djkP2SR2qhEdfL/pbQzgAtI
6XvjthGl3pH8PqBHpuP4ZF7ll3eutBHj2JKLUi7czcaf9AwQ4k00IQHRWyUe6qd0VrtY9E8WwyEV
KZDofyAPVxkrgIUj5PdUVvdzuLcKR02PJoovY2RGg2bAAtcqzzZt4O2WQ4ga33yHw1kMTwCUyvDu
EnM7jF4JVuBYAofa24rIMnbieFPwS3CSmcpZ5TfW/QGc7vdXC3Jw9cFuM77UDjTOORc0IFeFi6T6
zDVZbc8refC36aTXtwd/8F602+3VItovAwcmyoeODrZfWrWi48bTLGucmnU9VbqwTJ9i2wItsu6c
n9W37PGlgsC4jFsq2Pl7tRGqpoD+BlI2dUtklCU3ZowFwcVA6nl5G/beLND/yJs+ehnElJaDwDs9
hGRBfXf3E/YbQ0tbNMIYNbE7fZ2yJ675wkyICTOJlKwfhowZNr36bznGcv9rPTB6mmhxbtjujZ4f
tw6amd0MXCWdSYi1X2PiVNTDZAMZogLUmmob1ETnlunN5ug9pAtkFio4SE3WZ6EFzuB6mqKba6fz
msXnnYJFkRar0sKfrBstapxA90EuHd0r9wOfE7oOqj0Eto6yL12YKHyqF5SopoY0PQuix0TXwsCS
YZZaiUPkdL/UdX3WQ17EfDId8FCOh5LEw2lEYAFYWXzyJFmyfZdXqxzmwRl0kIWwaPkg7ffe7xvI
h+fNx9Bzb/ndZN1dxL/2wNn3hsXvnZEMwXV5pPb3mV5sFj7cYyqz5NZC1Vr6E+s+dJO9CIkRFWj6
ykIu+YA4WTwhcx2f5DV4ABUyHFmkVdQM5ZvYIvh4OReVFP4o/e1x4qjhjshv6F2yoGZlgdz7irEF
3lj9t9/0JcSXD2Ay39NzP4AnpSYDsoBvsCAEGgdqSQ+6mT2HA20sUCZk7p7MBvFn4kKU0B5blyoZ
Ovki9CLaYnKQg69kNLARyNYCIrogWknrmqNFm10+3inmvM7vTRHf8roy5ZOgwFPebHc4iA9DjFh0
BuADU7psk/N+7bRdgKwrG2DhEc70oDtGEF/uSwv22atGApAHyQcU4ClQp4yCt9hD8gP9mr/XB2sp
Ol37eW+ZlggzC5mq8kGsRBz6lbOWmzxoJ/1iBcr85ZSNyAIa/Dq5XQDbGXC7uv/h7Tr8mfbqbi7a
r3WuvgBWPnmvnUbrVKQ5uCWfjqwL75aA4zoSY9/sHLo3yfTDekYpJSjU4VKpdvSmtwCCicPzgXN1
X0rx0ydhsQt5d6DVOsnp24jxeN9taa800fYMfa+CxxpXjLR9K00YPseb8HHS1dRgkNx7szOhRQeN
RscdZNof/m+Gfi1ITQW2owx2ksityeDIuGexPQCFZmTDXDyLUCqY1mlHhaWOcIRGTzXgOBA5KopZ
YgP1/KAunQapMsCDsiBDnb3QxqcWZD71E1P4PdCzb/xsvwNtdIk9L45gXBgTO6s6Y3g/YH4OVth/
c341Ckj2+1MSwD9i3ZaSt0rDwAMTmUSZDjxCbSXhC64KuJnSBQeJE14440oK/p+uCTkjMjwmQkaI
X/FO9mHr02qDojjKlPOUWg4ORcYLVi6V75i02M3p8SBajz2AAvw9pT1WC36ssgsP+N+ZkY4ZmheL
eF1OuNra1sjN9+fVre3QG6vCsJ6jZRWfHM1CFOwiuyYGlxvGe8oD7uCwrJLj3IzSrNjPoEtdwMHr
Zper1t1glA94qjhqOrYYVPyS85CKqWZG2DEHF1C39MOYXTivZcHqmJntK/Sr0akRWCNBp70VOrdK
9AQ/Y0RAAbUv3Dng0NxGEtaXBEZL8Wj0ODuVAB5pgSIW3d0SOViME7ju+kTOvgVtVxZ27u+MTtdw
JMXZ/4lCxb3WbtGgRTd9DujTPfipmsPq181GTDPruQ5xCV17081OZXmK5JHXGPZtlMo2JsRxgn1S
xe5/wcn33xqhswcz9gdo5KTNF4GylCZ058UQ4FUfBs0LlxB4cRZmdk146vjIjrcYM53nUIVDx0LP
D0C6+6amxj7VT77EYz+3yRpwaJo1hgM1jM9Yrks6jbw5VyozvX8kV7XTZoaVDrzpz5iSfz7NlFju
/RFYmmINuef6i2+Xq7jAvKiRrTXaIXkZ8Gk48RC9Hxwd4fMUHGFgUASZi9P8Yz3kjLrn0EEsgqOK
bm8UmPiLtGvr9HrtXF94vq9nIqOICzpbeNLySYxBsLmRs74IdiHVB5EYvIulmB53Hn6yJGZ4xPsu
7/RlnyiF8MFNpCE42PsG/+IvXxgMvHSTfHoxkIzgbSZkPfaV+O/jxmFHK7kMHMgwPIF8hRfyD76m
NrOmZkBlnjUEH0rWKFdcKToHsuFEDwr9FWYxPXM7TYTmBvJGqu8pypPQyW0kpLrVqK9Mw7i4cuVF
LPrOH0C+MBWHldGttZ+q7HNrQh3fI6kq71MM+/J2vUi30qd+05mmsZFDjT5M9VAACgfkF9Js3eiL
ybzBY6MWDI/A1PkVL/lAF/td+8lG1jNFa9H3XMlPOkV1N9QGs2kTfg68CAaOuQbfjtrSpvnj5f4D
SxQbrG+TRaoKbNL9luq95DpllLrLdMiamAjXfgZJ0tmbIKLcFmglmdqPRd8alp+S0IhjknZ8aSXH
1wQRhUtpG6h91WsicylYC/Jv5WXQtFcFPCXZbHzjQNwce/2c+9r1elWxbkfU7Y9Ader/ev+rOiJF
SzjMBUC5PjpmIsReTIf5hFcRdI/p5+z+InCuxwP/HpKzUnH2eekTZIuYWgNjyc52rjeHgJ47m/OW
klFF65D3/tZL/aktopCTQeN2eNoPeOiyerdYqzzH20tF6UDUzObwBnyGEDywfbBvfyxAcR5jaLeq
9N7Y1bMqp5l27NgT3hWfILlRTGLA9q6YTXsIeLUmvFc+Kk+FkV3k3VfGhMEBv/PWP2IDyK1Gbbm2
W+1T42C26maqSpkyPQIiIO+i3apFHjorgqIbf9bEgj7JKtwpyWMu3lL4FAfOa3vqu/Janx7A7O5n
cqwZLhv3QoKOpWXnJa7TIST9F44FOcAipCi5rzPp790WBdQsdw69WBWwK1GGMnb1sRun7cGKTrFc
75lgd+g8TE8ae3PV2vMpoG5+EAe4XxLgMkPZNJ5mjcR+pu0wNqXgEzbnfFlh9nqdryC4kT8ZFPas
4aE7OW3l9cSUo2YEZVdWc9+tpXjL+9/fygvx9e7IYgSmqF1URYrqmBDrf4+6iK+/QMMu0+t44aZo
03XvixPe6s+Y7mTLx4SqQsWGQbWCoslw0GH/5rXQpnn5XlJmUrr/fIpqnujegrSyYdpVwHKI3m4D
UCSF4flzrwfMzJzxhBdY88etBf4NYOBJAT01x6bvuAnHJ7T7PhFKElSssZvhk7+kMKw+xiaeJAvy
KRZ8w2trrAJsNzIstSWJIVQ3tZ7JSOKLcFkwvFg8mXCKMedOmgOjacBdmdKp9Imqh4Q4RomNgipv
mGhYakKYspC6Z9YfnWlCMDNxMC+GWpOjoczfUbrStRhomouXDmLKZqqFsoo6dXQh1iAeVJ/zek6n
GS2foeOgRyEf9uAjGnm1uCPVQ8dllja8VXvJ1vhbz/r7At+LmKaGb2wEe5CE6jMZlcGWGwLkYOHQ
KvczbWrECwEOgpwodkXLk42fst0p30BjAvacwaojsk9/hUofysBMQE/LAxDCSB+hq2WMNrcuSPvq
cDA1NDQJy7N4SzT7qn/zUjqusiPP6u0APWzO7c+vuD4OjgrZuWU/DgxkkgEunDMr8z7ZfxDG98Wg
FYrUBoeh5M2rYdljKQGwAENZZsuGo13UDQKx42j9VPAaYRuMFRzBMiMGrYGYJFS+dGpBLLdJETGJ
8lNC4YuLbRoRVBEpiVEVaNY8ryKEnvQ3X4xFLTxaxrxPPFNtmwPfnYWVblm6URZZ4NrABr8QHbmg
XRfSF9zSWhXF7Warg69+GTDi0/ogc8g8TLuAmLBdft6ng/DeVnKiPQkkA/oGYjjvV+8KgqoSyX1v
yjXLWqKp4dnelQcDyP+qQ2wFpAQ5jt8dJ95mB2iilSgpjTSAFwW4In3VEMI4gmQXiXHEcKf6GnhW
SsYF3tf6WzyrmJ79OrFyx03++/Mq4uB1veV5pXCp8PjGBUeIUlOlI2qWtZI8GCaKtKZKf3jHs/B/
U1aYXwms3THU+ZfH93XQ56j8c9/de8cdkTx6/8NVbrykjSreOuWOhpC9F5eJUOYg1bOjoGxdUI6o
8BjUXjuPITV9ln33ffQ3DNz2kUPZRosm5DbTrHqFA0kxKYt+6QXeWl8yAazWgLUatV2NDKOr24OE
YLXds2AnSBi/8BZnsGDfjw40KNFVHhSvwVid4/AMgXxhHa5H4DOVl2fhGfMjmB7D+7fRp/mTfpJU
37D2HchzoSX5XkMGoZcmT2OY9iuESPHHtAe46dLTYM9wOD8tULYNbon0s5NcIDWpYyAMjpKymRLn
AhrXk0NISG8BCc9Lpub2XAH9mWYIZxK1fJp43VLdCh74/HpcdMJTfXGnV84qHiQ3Jz71czHHggnt
YIfsEouoGC0NWdLeFifhsOf5TOMYBRMxHGNBb2QP1KwPuyCcv7KtfORDtIcXXVJtMsRAf0g/m7A7
ECaZo3RL4qHu/QU3Yanv11fIi18iXNRayw9n8xEgNy+XyoKUYKr4NcoJUF2VOGhEfmmZgeFSBj3a
jGKYcHvIPgM92/uZNpNSPo9vC7icO4ckZnNtzpIDkQ3SPQPhkWw4qJ/TFT21eyjWyWBqLF/BXuoB
our7yOgEmguhf/9GqmMtkN4lpFWIQDESaTjx4NDGiOV+dQP+Gc1ZCUIYbNiTgBOBkYvOGihuySMY
KGFPHxmzkGjxmWACovwsQ4b5U8wMwMc/6WkCeAyQWTmnWcj1Ur0OqJ2JNkz9Ucvk9ElZUsFQ00I4
2Cl9vJlKGZuvV7N+eTjJ+2r20TLrzvphdoHXca4b/WlGtFygxBFYoBTC8BVJIFZmgTQenj5gc92S
gQ/wXtCJurLKT1ydhVUMH3Yj1WB/0TCvNWzr9DITlImM4JbFBtxG1lAX1T58pvLyu4+xeI3PDSl8
KFLzPAktaTekHrbG/6yyhWPAd1l7WCj889PJ925BxO4HWNrahtTizaxsNpfQ2rskU8cL2/LMywp8
rvSLiu5zYj8aq9qvy6zeiH7apujT69ArU2c0+Jx7Ilwp4X+omNNr8tO0gCjkyiAqdvHA8owdy+Z/
x0MyG6QiQ5qx+VIkJ8SfWb8G9Z2q/vL6bfr3ua6sPA6dhYgPRXye1y9gatzzQzlcFUEL863VulRo
C5zKeSUXPez9TGhooZmRfIw26aKQ/k4ZbHOcstnc7Vxo1zkvp0CfVZGk+8xG8SxBeoV3JPh5vSm/
3wh3YZkfNqc0tEKCYk6yVfY8w0PrzNAfOpStpdhmIJRSVOXdxNN3R+7ztya+DF9mwa167vFnIxGQ
e/XXYmy3dIa+4rSgFC842VFb1IKRimUMcCEXAjWV56unwNmUfyoQ/ly+QWbDksc11cntee0J4dIu
hTsmBjsMlztK1yI2JpIqVPomHg1qvOyXJd5xZE1A9fu70AMaUcn6PgATyeu+T6RKVU0PMM3nXxyy
zrFP9yy/Z7/FoWULBrQX2aE6vpEp/F0/+eO3pZ4d8Klltt7lfkIFiDoJHs5Q5/dx/SSJV2o/fte0
P9wRCSMcJDoJhfVpH8GanVt3Q5XY8n3kezrfe8egoggg1/OMcKEeMDqvDSS0ciBeGXy42NBIHpb+
9K1DusaLmnQW1WPPk+Cgi3ElC5tOy81oUhQUf/PFQ6MANyjr2PkkR86ZGT2UB7N1EbN/Zhz4wdkO
77ALbF213O2+uk58TomkRONO5t7KMA1O3eeaKshzOwkNXaiG5gQcFUQhH8lPz/q4V+8LiLHcCxQE
dAwRgtVDAEhX6/KIqvdCx5ghn9i5stxxZM6vCNCb68GhxLc7t0d5hbNMZHMc0/MepN2N4CBj4MYk
fUUmY1zZhPqkTLJQd/cfA+0DdVk4siVs4FNJ4DYk2ik1EFb3BOlMPh/3X2Jl+cNL5ehVbX85RjCr
N90ecHU3AJKO5S9CsKzk1qFxQxdd2j4Jnx5W24TuZ6HR6M4v1jycCVf/L/6WZUICIxNDZYEFH4gJ
ARTGfu0vClYPYzXx/ib52Y6/NHUMXwEXfKOjvRhZKk/dzAMuuE6jxdi9PYg2unjJuEDobyxnuysZ
gpa17eBf+JVrAf/mb5MSjWPnjXTLRJ88xY3QuAdQnQ6A2QEg/dVBEdxw/tOzu8nSZRPInwkLct0X
HHjelotXnuFVBQ8UxRrJjkrO9NS/js5kqF8ojICJzUAhVHo+1a8VMByBQdAhd3zxXvZhaB+SbdoG
3oPZJOsvW22r9xBOxulQvESd4Rpi86hUAWDZ7OWww/V9F6e3yx/Y4PbbPJI/0rxRgmrGHlVFRinb
M67zTS54ATXnZRNqFLt8mqDDK3Y/Abl3YHk/PhV3HZ+a04WPHYNW0VSXj1Dm8qDqkb+FrmVMX2pc
Q5MlFVD1aArBA4IAngHei2RK6OaD6yvQQ3wK8wwdsjwcKoSL4AYOF8PdVD9CNa8w7NcgChuJl+DW
7pj2X81nVdWfIVewcw6xdFF7FF4O2cOBAvF15j8CBz0MunlVbrJYmZwe4vPpJpdGItp4iYT2bsJP
tx0vhwnI1CMwtKMUUJ2pfZmwWdSBp9r4eLnJIzcvI77wZWNgyo9Xi6Ia18JZGkiQlAq9k1+6O6Fu
69CyBnNrTA0LXEtOU7sqk0JQhsPGTZTtMbhfQKYUJ1JGg1jMoExnRt3tIk9gTa/UT3FSpBA8AhZe
OBJnfhnisx6FZIjZf1bVBoYBwXT21kEEL3CC9STr1dcnjH4CGXQmTKrRcGnNaeWLaTO6hfjcMUuT
Y0Wg3bVg4cknnTH3nWQCsOKiHJSna1QTjzSIEfKjax4Q7skxZucQVw9uk1g/7uhDj0XdA4CMpxPk
vOG4i0sVFr3M4Xuun17A3KlhqY8FCz2IICrxjkrzOsofZITQ0t0Kx0uxyVn6b0vt2DnqVodY4YV8
Z+ZzN6Ir/kKk5017bhTs8V93Ux1fO5qHoW/6LixP9RJfn9CvAMCrDB8i3BgK2ySDz8el9gAYufJA
yY16a6iX8WzSa3vt5ksY6QxgbqSLUf2HiKaYGtrz6mxLDbJFdhI7CD3jq2/Gsr95ck9xbf177wOT
VOBOmDY34YbF7Mk7osxeqJVK1muh0XfPyOxleOxf7kn5hx2LuiBPyzG0opIJ8bGMZccG5cFWxnnh
XqUeTduAQgUZy9BRjTTNRxHICMSFXS2Zlcvt0duE+FZo7ajPu+91sH+ALPUXIVE2n5bpHbDmPbqH
92SL8i9tMlZijiB+78Ud7yVgWOOywOdEZMgha+hxHqODZm9MnQZ6bp4zyacbwzMk9cxWBwKoy3LZ
v/NTpb0RHMCfo1sEOnb8JNbF5IVtYkl7YnjyYVZMVZ6m24PpTvOTWiD9/F2xBLon/mDKGdl2oi5K
J+BmuhWGhodqvqPZFpH1Lkh1ch8BENfHnTpSDf/engZxJwqy3/p0iQFOToJD8IgqYVV4qnsQIEUB
QlmUrOozs7FltJfW7c6A+UDfcBxXp4gBqu8Lio9ZNNSunu/nE/0nOk6mVuGKZD4S2qcWwn0RMtKU
K7V/NTZXVUhe1gOe8GNEluhI0w+MMkHnxNEIByEoxwasQMy5c2SjuK6uAyB+eFk6MMLcFV5bUBCW
HPii377Pzy4aHq3lBVcMPY3B+k2jx0SCmNjlZ42drMegtFz8rSpXwyL1wwMEm9Muelij3xFi5lXN
VOU9PW6/9gW7YcndR9w5yF3C8XTxpjAql7G+BADX+edjpzQlYk7UHScrS4zknCW/Zu1fV7ZVspJ7
7TWtwWUJ4YZouKJoRns9qIPJU1faPpDI6q5gtIg+R8r6kM7U/s7hk1hCXO7URpWvZfE7JTCL26jN
EbLPxLDqMy3yQ0HjcRja6I10o0BTIe4uQPztDHcR3MYFFa//bppiyc1BYTogpMIkqIoeGvfLCek2
qSvDF5TG52BUxJCaM3M2FEUEt9RrvuzOnIATNAlPP7YB1FsuCmhxeCv9DWGhd/ogHNE6T6L4H98J
HV518c1QrV3fauNnhUQt4t+ACePCeKgk+8SKmemSAP39w19saTt7kgCN4UvFZDVjK67BbQn/6k0p
gfrydif0zfPhaHXTJ4hEa+QwfK9+9A2T71l/LMS0LT53t79wMESi+NnV4R6u/g4agsA5SFaUnYfP
/TiCIKOo3wIM54HRkGvSwjOroQddEnoY7qgMNXr8wW/J9sz6RjynS23Y6eDdJWX118qdl9/QgWZn
FuF94mNRllFgEu7hQjLOyBeUsJCWfYAd9tD2x64EZtRRd1zHQsY8LEtFs6ezio6SPY+0eHKh5OcI
ZI0+U5Iusyg5dqahFBnXIy9W5/HCXyrRCDk/X5mJ9VmAOBCkUygr0JTAqByIOflfmpAutOk3MH1T
Sj3xT81SItNnZQfUf7l/gfB60e/+ysG2RvGvcX45/YT4xud3oQN1VdPWbrmrO0X9ocx5mxBdkXuZ
XEMv8FoQ+a6IfiNgC0UaHfFhiKnPCJuNl3qA5DW270Yk0TlTjDZEpAs4aGxh+TNiNLdY93lPenBG
nc9U9kNEE37uHHQjTDDA38sPTyH+9M/+OXohD1YWSErdQpvC80BFFe76wbqtqfiAQj/EXU5lcub+
Sl21UFC0bMg76DTjVHdseDahT+uRvIehB6HSDcRWubipjNImcUXV8O/cTYfo/fJyRjRcodq1hnZB
h23TPE3h35Lku05HXsuxTwkO6cHl1qX3tEl8DtLEV5yaF8i3i06A0WP5Il9tQKtSK1LCinicN04a
8lT0HxsiT7FHSHY0sjelX268XdT74cZRtYYRUE/839kD1DqdNgclSO+hI08TNdKjFF9gSkYRbjew
gY1as/2A0E8TQKUBvkr3yHdPLEgCacxWGw7gXizhs/CKF4hrmXynIJSmM4FKqty9GzB6qIr3Y4ub
guG0KEB3v3GMW8IcVSwUx2xNadePOqC5LfoDxI6qVLQUCNr1Gjd98sRrZXxhXfCOiS+zbehrLcoe
RWnnvsu5Tx9I2bFrRVhW13wAFCxa4HmvhEW5se7jDRnYXpLHhLFKZd4IFuuIAZwLVTmt07jtDckL
iU3mNJBUEn6tXC9Im5LsNgivAeZhIYtoHPpy7UnGB7vUyAhTCs7Do8lXNjno1L9UR+Ct9matVhgF
gWA04cZsND9cwB7NqOvFJ5VTGNEEsO5f35bkdSD8plpWRWrTzQgk9BH+gfFcvDmgiemuE6HX//13
Srf+GwO0T7Piqx1mIA0Lqfx0nL6GW+Jx+YBVD2KU+HnsL9GmD2dCrGx8LnQeDLc4V4Lvdx00WVSF
haWSQhd3aCml7DyG1xtUjUJwBTI5jxe2W8K6S/A8+3+D9fjXFXgCuuFIxdXHwx5wGVhTn/FBjQYo
k9boGP23KZ2frn//vAg5hDxrUpUtPXkpZnrBEJG2CHcTXpHhgCp8FaD/bfe2khGrmxfMEjglKyf2
o3hWgeRiI65CU0oTL/dAw6kNAxyCy9T5BkbcsO926ZWsA5kXKp2UCEEQ2Ywjk8c6PpSzhQmfqWbY
+wwnDJFVpWo9+oPD4Zhf8kaicbw4o5wno7IfPUMticg3nzRoCkslmctOCaqSKbr6XrQk+C6AlCW5
yI0631Wx1mhNeVcVLEi9fEPmCKN1soTvA6/8gfThjiw77HhztppswpFjT4zgxceqtvPk3DuODxRL
7kFVyIAQvo6il2vnptSpJCAhqijPehkwLsBW56l5BZK1SGR+FWK3dTikqTAt+Lu3kcrP48OKlaqX
v3v/yQI0/mt6NjPsx2xc3UUz/8pWciAb2G/jKuEgvrTz1zwEXpxeZ60hqaBQERX0rOla2ut8cCbU
STXkSM68mPU0myHtxJBUznDEe3Mxe+ctFoKmrVoPidd9kJ2tAYO4TFqzbbdNOeI9nOtIEh1HAP9Z
6ls7uMbM6sc4e0Z52LzDj8HXYpupbVkCKbyOO3mKJbUZSdBkcLtpUY/6uckMcar6EpPvpBWGZSqR
A4S2J9twiLXFGTjarWw/DjBmC2QmyBuBUoS7tYXwbTtz0FeOxxSoW+OE7fifuhok33db6JLiZTLr
WG26Ai089Ozzs+WjE92+9O4Xg1xePg71Pe5b9JaTGSUqiTdD/AUK39wIlG63cTEkIqT9ayW0A2gC
QczTcu3yl1RyrhehZEAxDFWCSxb4xIVpoI97xULXRG7Hlxf5jVkPozqgbbZMuUJBlshlSCCVZ5TA
1HQLaQEl8jWYQiFi81las73Sf4hlOgvCA0YZUXgKv1mteurtMHOdz/4sxliYTh7bdDL2iqpxjO1J
VTKDzi0AWrMqAsbrEbecbYHRFxi3UaFfZ7N5+NYuBBIsLd0jat/ABKWwaETpxnDJr/sWP0ISIbxX
z5Fh7N2peHrPPE9Dw33fHI5PvR0IfEoQz5MYp3Uz4kEpROi9dLDb/PKuuJC1zI3zry/5SdDuIyS3
gQrDCNzm6Y54BK3xLYZNnSuzAEgWbLu0/TogJOgWiNOhr+N4YRUFakuEz8dI0L5IhZM7K/Y7MXlF
aisa2UpECH9D6CSMDh6UfvKIfVNJiyHq5zVO7Chrl1QHh1PF5R77VnS0j2KHaa/JnCoZG5OJ4x8D
P/hRP4DixQ4aQT2llp4Ts77RC/OubgLC3THcCXAVzGndaipE5A5QjJuzSHy6DYH1yH+lWFfxTwy9
9KOMsjSGha/xaIKtJRU83uJwMW0NmB2nMjUgrT5MEFFwNaO+kDEkcNxZz1AW3WA8N8/NQxr8nZxg
v9wu7EYEJZBvYt9EAuApyb+ufMM+33Gaxt25NubgUayVmJGpx6GkXs0lWtOFAyZxM/mHZGq+Hb5S
d9us7WCpCUEFxDUmvmSA9Ta/USIrfwAHtH0/gZ/Q8eyhMQK80zV50F74rgSG5Gby3r3bfM31kg6l
XZZcis+lOm8TmLTCbMGilT622jYQeDe1+/sQUuWrWIPubED3+OWU7t4TbLHx0QRpe1R4A15JpcYT
DNArqn503S/7xO/l/HGfpoYlXbRBYsyNw2G8QRJ8ERsZEMd6rxoUICSUyy4InP83g8I4XNR0CC4m
kaPWkWqHW5779/Yt/VLRl4CdzhZuPSrnffp6ITuy2IaPyga4RKxyBxFtFiOMBo+YVAcTdfbI3R65
A1tUCS1ej3kWSeiyPwAA7reCTu1ir6hrxQufovF207AHY3kBod3dXrl9mqdB6Oij6g9BA75v4N8/
Yc0NG59oySfPqVS5l6qz/7H+D/+DyqF5xleyM5mXaCurEVK0Byvns6BLLDgX75PbD/B9pDHzw5vX
af6mFv5R0z+PCzGU/kW9JLE4q32xo1qdfvE04QO+I1F10AxJInPP/mg8Sr8cE76lj/FuzxUe7UTi
t+CGiNbNgSYll70tVKdxXBnYTmk8w2eO4gPLUO3fim+PUaVmOiAD1db6r/0DaYL8UtKG7G58nxth
qAy2AwrV8gjJJGZcTFrDZawJvwfBP6l/UXZTaiBVAkvKpIMjKaKBLi42r2Fl1WKnFvK2nN5KfknL
aQOSP3qryRv95jLJmLZIqe4FoD64Q5EkesXKQWrgu/pTZBeipgFRgel7d6BbS8IfkdLC20EOu4ra
RXCF0wWyloPy14k4f3XztMGiNuf81PXsw2wkHMfWn0Vd0DF/8pVrWn3MsYzzQGq2MCUCi30mubVb
N4AQwHAqaE7ZprA4ZO5btK3vY1JM6tTekiN2jkKS6meVF2+7qyz+YyH70z9qodro8WIVYB39qZ5U
glRyMcXjvDnaCQHOpFtqAJg0wcu7wdTUmeq6le9/x6YgSCWNL83ZPCutgi8RTJTlxJkyf3jgPj+H
n74bT6EdVJI621q2zL+5DiPgsMHf1I+dA3HmkpeX+fJTWsIT7LTSW68wF1Yg8VHhU/2uj8afck2E
BMMlXHLB/H43ewiDq5lDui4uiaDINAWIaV1PUgcMBLaF8cVXeHfwAJBvaZiELtpToIiOPYKNOAID
5tkg7jhNSSjJrgAZNiHNjX/nccE8yGHZzr6wMUZ+wcqBaQf6gyNLdchoh+c8TE2ybqw4L6adcco+
SKWR4iYrWJBcpjnU18d3EhTt1AjrmrHVwaQTLAwIBhrrSME/0SdCoseAT54HoXRrMHtMw98Titsz
5n6L4hrjYSZG3kC93Z2M+7hGGFhU2FfzxxGJgRnRnEKcsFEesgn/nVUSH8LO5ab+Vn7TrYPxlOlJ
zTLvHqZyA0O6NWuhMtXRxC1j8ZBlL7Y+euOaCQRVmaZ5qeZFueH04Ph8yO4bRA/noJru54Cw/84L
DaOu9NO2Hm7o6FlI/Kw5692eO0ddddpr4rwqjWyzDrfbAvrrSM3XBlM1STU/uy5cP8B/8HM77Y3r
UCPBmADe5k6U5F8Uxk/DsomueJYl0szC00t406bX5uVfSx1BVQLnN5WhpH3BRhoadr82lTu+jH7b
oDMQOSVFj+nTqyagr52+wP2UevWiXigIU1DAdEDjqPbY4fM48p8nP82H4BXoP0sQVuq3yKqI7AbQ
A7qJObHJ0bxBoq6WOPtLpHK1CDwMLpR0cRziwakLlnf2h4FRLwRhYydruotVmItnwn4CaUaY9EJC
xFu1H1/ev67qqPPoCMsFZ/VR+ekJ7nTqscVdpDuns4HE5uP7HNcjP+/e7IUv6jJ5g+PkdczRMkAU
ZfHcnbU7uKWh8JacFAIb6+rZbM9aYXQA/NxAt2xqlFLimpMYwMfn2G1wubE14dpVme+jbuymTnfB
iUvVBCX7Q9NX69zLd8vzLGJRXFbVIoOuXoEebaDzuZzKyLaGx3Hc005CCIHFjZO11miY2j9+X4Xb
VDY5nwnp+KJ/VhcY7tXHVcHmYpmbO/FFWpjQlecRVpsWHtH5wa26Xogzu+dZOWfP38eff8w3Mgd/
F2Vih6xS1ZjFbXIZXHnluQ5WXbqlj8rIqfqvS8ISE4AaxsM2HaHC9qSDzlPLRGkHxgWm4GFSArVo
HpBV48mQ+aPmI9YiJVxr+plnrQKKoEhj0Z5X0qrVH9sIrjLL8jYAQx7Ycs5sIQJC6CL1X3ZYv9Jf
ldBnqGWvf/LXSvUehuoO+V6HU8rUSZFu9a1xYMda3Kx2saqaDYuYF/p4oM2l/WBaxaOai8S+w7xJ
CPRie9jeCC24Jz2hyktcXfqvai/6iG9zs9UI52LtVMqZvo/Xuly/VhF4G8taW6biaU3LnoZUb+5K
weWvwoX9lkb17XohHIzdR1aJkyQXIIlFhj94JVdY8zBEFnKr4vBSxKT1tdurQNogV+Ul3Q9fcW2O
AmiZsomhuozIBn8dc6+de5UAxJxL4ZMWL2tDDxjXaV00uGDPBJzM0MuTM7UPkYj46WKccym35Ald
ilfFU8Bv2gLVnSTaaedOgGZzbNZDEOvhM9lc4NNIpRP56nP4DL+Ygf9Kp36JXq8zCevHRN0SYRiI
VyLY/+P5dFU6GVjCxYR/r08PEgbbudGFJJHdPexMK2jguaflQ2Dt/YGgSRE5YaaiJ9Ov7MgX1IZQ
I6Yg1kPe+Lqkli0yiygw+Fvi9mvTfazKA3kxI3D6NOWNVj+3jce0U6vuHswgWRw8h8T8S2V24AFt
6wFoChiFYEqhsxHXozhBIX9Qnk5CpqNEt58BaoKlZYjgw2Pi5bkdSIGtE+ZmAHGKRsWw24i+Gd0c
8QXkgpRN1LRltVeu3Cm4pXy7l+/HGQesnPAEDDismbnKLYu2mrXIHN4mDySyCWPguRTKmYGLHkBw
fgOJ5mhg7yGc+84IRszoY+t7Rbn2LsJGOcD58G28yW4qky/5d3vFAyT2+odtSz+WLsTxd9I2nkeL
Zm8Fg8j9RjP1PnI+uqWEFGYeh51sWkBoU7AteuvkDGC3uvEJmXojhC7hCTABjofB3D+S/xLtRrjX
zPdBkKwHb+TSi32fhb5NZ8vgV+sZoj49xA3lcYNqdkuFHXGVdzv7QZVXbNNhrHhORKwmuw0k/Ga6
87Gfv675GOmHU2bMkI/w4BeY7ewVhUvU6kEgUMgjJOBpNSNS4ha4EScUycLLPpQUDgjQ/ob0rr25
pY9HevAQI7aDkNVZrqOb68rcD1zQ/CzcD4TxeJI1A7e0js74a2c7Qcs31FokowoTaQ85GYkq+Hfj
9W3eqmzoBfFKYx7Rrikb2L+kw0GQaQ9zn3Ie9ZSFgPWtitPK86DcW3I4+BmX32m0NtC8LUzzBGBD
CAwBq1b7Tfl56IxR44d4KZLNJqOQ2nDu1Zgd0gPZefa1etVyKZgNUDn1dks4vsncP0cR7Ug50UJk
gSkP0zOYfxsGb7/EG6NpZ6WU7zj5kirwGivRVgjcQTyeOvm/A+s7o1PBfvWJYaxDQlGudaLegdF0
taHXdAX28cKgwBZYnm3N4B235zRgg5m3M4Z1T7SX8ShGjMvU2Lj9G9qAVsnnQjxZ5o/EuwOTtPF0
fl/FTnqzl6rXwF3gFIM7mnIi0A/RVtr6J1+ov9BVGGmZmd14b7iAflItjSaC6kbkNnzxUWb4zf2V
/tiY45KdNYurblsSrULpofd3Ol46JDONOIP2BHdo56Nz/6IwdikQL27rSEf349zaxbXs2FXDH2X3
G4aYICAvF5PCaw54bg5FKGZshGJWAX3b3Rn0DXIY/J7eEscUcZ6fe2i/Y/QTIWo0gTofppjUUb9I
0Ms3LMgps7ybVDOre38UkhN0utHbbfSmseLv6LJqBkxHpOqsW/QEV4XLXkjrLsmmoHdC12tyBJzi
oiWmcajC8pP56KE9/iHXq4cXUpqo/p9xFDqruWjU5pvCrODKMIspn+RVSicg+g85IvKNqgwLkq1M
ms2q3AtroaXQuK46P+z3rfkE4I1xgejT0YoMG5dtgDPJCBnH0lIBQpF1BnUQTq8JJhvaT8E5Q6xn
J3EJRIDJbPRwlTb80UTu9vQhPUI0iKaAoweIc2ROg52XlPLThaxJyiYJ0JDeJ6Nx8I1YKOalYlp3
c1aEGx3eeOrpDAjhvjni2pCqJuumCX/c4GoSEMWSf6hYYGfWU0QpBaZiRrBSGmI2amU06DiggBpm
ii+zfqqVYKWrA9Z/IjqIYxq3RU8KG1O2PacG9rVSKhhZM3YoXmoquxeav3mFJFpb8vZ1L1OShTC/
CyUZil1O9iaRvsC/OQIB/tDlkEiap/weRdbJznsb0SZvNcPrDrQAR9gX5PSrwwZ/V6X4WELCeABA
70dM9lI3bLBd4QxRUkJ9dsKjwKYCQd2S8SdFg1r2XWMvKLHROghgrQVlhpqgef3iUYLAX+PjVjin
fWuPWNzpTH+8UvVruH+ACF0QLd1hcPrJ2+Tt1ZND+F2zLJp1FcGaThXW7MHp9DrZlnrHoGfDUZiT
PnsBKL6baYGKG4uPsnMRkY2vko/jcQ8BS0US2BAT0cWsiZNc+OakVgt725+EdK+NRcQRZWu54jkS
U3gCO3iijgUi2AaSy5YSU7cYoVgt3VhPTdTGiGSLSkgyFQXoaUh73DF94T7qRl1gTvFBjbJ+ojyZ
C6uiHzQRwQ/fsGNgA8trpIJATO+2hqY+S6GbeO6mskKQN/SEGqwuS9QY7+INy6IOd6CH/GS7kU9R
1q9VIEJ/vHd9wfP987gzdwMR7tuZy2QK+R+gS7lNJNTFk8i1c9WiJ+miAgJWiJbK5EKZWcUVQ5Xh
g2+bpbcG9KElFb7j4t0H49+4iBTwfwb7lZzvyIJkZgzbfq9bif8mrLcAHsrXgYA++IfrOCJE/QZW
MV1YnmGwetgKUV9Q6zkUdktSkt4sHvwLtRER0bhGBF3RB2UrXOjemfQv96i4QSh/j761KE9mvoc+
WFUliSkzIXutGQtcaPVre1Ado70+96JwMf1eOJly0DMojy0U2sjYNDBnaTnbWmmPWi/9wNlxc47k
fEhofiblEO3fRoUk/vfKccClhNlnaNck+hHYcw29NJpmdK7TTCQONHqGTi2yZbBvehEDKtVtq1h0
5HivS8cmOUbqzpVuQ81FD8GpEODDNajLw1KUQGh/i1YHjd6kBW9cPhyJeYwqgSNFu6CoJ+yB+RJV
xUhm+F1SsEQ7iVVyGc1vOc4/CinVi7Y8BQAx+q4wOcrx7a6GYQ4Snrr2jpOSqNdNlKVGmt0AeH/g
5oQR4j9v0Dg0gKH7iImu6F1nWTav8oxy2sJKbj5UN/9/x0Tn8neFlVGWjtRGmQRJCFhfL3C2owzL
MqnUBOQigrBx6bx/pn85MkKpOAyWDFptdBFD3vsErshyyUFWDxooOk+EW+o0QID8urkUntlN7gVq
9Rd5mePF4uPVoO0znHQkuTlwhyOGBfOR0D7LCv5hzWyD8bAusedwm7XAtprxpycftSpFeFdu+o4u
VVg0niC8HqzIkjxn0LD6Q5nM+giNhOjewjRPzbk8Jkej7j2CsLoING12XHjBIuJe9p5xuhKImWj7
tIqvfkg6V6303rGvRHnxBCjppSOwQ38sYXG9JWXDqrqCARS+uVCjz4TckuGBv+cKNJAVyYDBImUM
PJz2QAhHt+Mbaw0awwcVI5o4fx57Yu88ti/EzD5fUW5fgZ34qQ+qqESZY5+RWQUyG8L3XrfqQTWi
7Ptwi+0cpVhsIcfj73/F+uVwHDaZCWbwnC/z6iLlfNheNegEMF+9yF0g/U/gGGJk9K7rP8BWhrDR
OKHVXdBd1JwXtx7zpY3Hf4HccZ1G+qwKP9AaOeclcQGi6WGybQk+EZwMild/+O9kDbVcPjRHZmdI
/naXcrmsrICQoYiGmxgPZcn2qjXzwcHrWwC/UUdTcAXFK9DxNPgW2VSXbAwPsHngWBjmtYp4hcW8
d/Byu+hjEP9tkvsg8S1xeWLDUiELbZUonliYtPcBLSf9Do35443bJUgMFEPU9Pzao2PKypimWJiQ
y9t+oN4Ih4g9/6SHsHTs3EaqjEOSOImWFKoEG6BQFXiYzNIafoxbZWuA+j6YwHlEVTXdOeaUyWSh
cZxFAAw9YSglxhXlQpoGWpI9QodeG732fWNCt0YO8gXwcl1xs/RD4HS4jdFZayqS3KQh6ie068gu
24hM9PzxuLnKJMHS8J0C5+QY60jOt8U299NYnSeDo479G91lUsOyMf9rn6AvSO0nw2xTbh3jFDgN
Saz05+A9FyF1XQ5IPHoE7j/YTgmrU3TlstL9kWR9ywM75ds3jLUT+SUuFhh5fqSwsF+e2xURtrUB
ExXjivxds2rcHHVYjtv8FLStf5bch5d/Lfc1KCCYfuRQJK0egrJTVCkyeJQ2C8h0dMNC747vW5mF
4ik2hCY0FmbPqW/eFClsLlbVGf2z0ZfWHY8guHn63+6SMj406h5n/vyzgrL4+SC3FTWz5ffGJeqq
jORw/CWEQbdoTYt1vxRCC4LSnDm3AFlDcRLkYQMDfWAergHW0v/belVTLOMCDcw5rya3yYCD/L1e
OjyogLA9q84I95DpLPAf20pIf/F2E5KIRiSvELkX/9AhqyxhFCXvvY2bxGDbFdGYsJqE/1A0XwFJ
5CiSD6Qo4H/JNI4LsOO0XQMk2syOL42ZXYdeytV7W2CEU6jdyzYEdlg7aYCz0ZHaF9FBgLiG/hRp
zgw/KtLhgJ8nLFoeuJftdMZOvqXKQ7DSBSFoCSwJ6JXpr5LSPz7VKHZphIpCHJL0Z6y7xAPAkOTU
dZOarwhbZT8/43JMAcqSWqv6I4SrEdG38pqc5Licqwx6XW0JTTR2YSxYBxZMexaUx45Ho6j3Tl6Q
ULjI+ANkv0QJfpjNsUBs6zyACpjf6lEkzOwV7WEAPnLq07ow3I0jjp9cTkT2DAZsyhzEZYsA4bSU
qGzJ+Qc8XudJByoHY5uZT8P0FuHs3AMGkEewD2XeHDWqLsUahcCONgRwZxfSeZK5j4SlJRnfsC/Q
W3qTyeIH19ZHvKnv+Vcmz45FggBiEiOtjymyS+unBmJ98rkdwM3kfpdtYRziBb6hGdug+kTs2p+Y
CaFQnOQOo1v68vJmR1YopK6hafgN9xZ+aUu/sLfWR4K2rYk/tpUy09XK7KUJcpSyHvpGBXvf4/WX
1TYU80Ueg+AR+01qAi0K/Yd/MTi7BjpgbyjbTxqMhnwc9veLdB4Z3DhZc1augBj+MCVQpNsSAnor
bdF/+FZ5ZZZVTlS4N3Gvw7lVKDCfFpCgVC01M48KQTSQE68dFT5xI4QYfPHLxzSPsWgDEw2TnwjP
FpA8pkydo4Tr9F/tgmWe2gqocpX3hyMXq0SwYTdzbMJtrOUID/CRzdesAcNkLlSwYwyuiHjkefsG
MZ7E74QSwPXSj9ylPwdVpNWSQihRtak78OM3CNKT8J5FOr5+k/HP/jkM5aQSzvX4khDubE3g1TWY
0hId43uLNShOMcwi+sSXPzINN72NV65847ouNIk0oXERXn+bRyOAsPOSQOKGzzG346ouXz9Sdtc0
yypEKVT0zSrq8U6WH/Az66K0RY9Cqm8ABVCCKe2pLV0TWYFOgUsQl8fOtwAsdfFwFF5pJNDP4lr0
H4O7PjYlulh5CBtDN2fiCKjVcgkB8eyUm4k3dXN4kLNtVgv+1+Rl8+Z4wfogpI75RRWOWDk6lbVo
uyitwkr+HB8n4IYtFwAj9+lYwbnYVEPfihN+2Adys3VDegZjBzmcJ6UoyuJB5tHyNnA50PACGlz8
4NGie0wRrF4vc84RlRywwkw9TZhoprpLeryK5E2Y0wv1dUXlvA+iPyadebjyZLcLywPZs9L4plii
8Lq3i40nrA6bn60hKS6zyOSaw+iKjpmx68laKaQrES6r/0sK7KZopeL3lgCS89O1qPbdWm2qILCF
DK4O7rhBwuJHtHPi7FaV/7/lUtjvcFCxOtA2w1jxLhkXdTLl8tiG87HifT6/5OzWxGwZBmPRjydM
lA6MUJ+lx3xljkxO4Qv2T8gohAmgLuQaIK6nLGrzjfqHux3T4KIo23HErdHCw5fvJvzCOLcPQVDO
hgzMXyANMo2miyPhmOUW8z8POFHMk9YzARsK73WhxBGU+w5vvkS55RJg0ad7sUo7akipYOGlvNuS
MFaMwgS92LH8thDApsk+Bpbf5gG/sQJy5D6XDujpOTfiGkFX2z4lLtn3XBXzy4Yw+CZNDbnqTXiB
WGf6GSvBmKT8/qMsqIoFBuJNxLSrsz6XYpXMEMKuf8GiMPIwbnnVQQz7btqIgOLZj5JeTTzHO6hw
aLmY0NLFuDXKn8K6ciDzwvTCZ95a5yNSejCeBKytX0OjLBosOdmgP9PNCkH1aWNgJ1CVPS0gaqoU
ula2YZXyvspJJuUbu8xlLAGblvjMHPnlyA8vN1abVPGvUHOZ0leOPYoHxGTQpIZWfQ8wEiLML82L
D6uI53TN+IePtuibksHHPggF2J/N/npNkw+klILUDwBKyVEjmK1LDg4kgMu1y1hdT71a8S7u/mQA
vtx2sAxzaSc3xJZPU1XlbTPILp0QmkvKfRSYRxXko8SitGziCj3RpODH/XNj1yOyZSsMkYqgVrY/
fWjkRF5lTNA8U4LT840wFLkyXVDZ7WBSd/T7u/BsujTRcccKMSGLP5UpygWip4RzDwvkMgEiepVq
siLz82ByLMqrvQwRJ/oM2aAnSE+I0CWzZgmlCzUKBT0sDXSz75O0y6MvcpCtd2OmaYqunJzcB3FT
FCH8Ezd7lrsmkHhdSei3OLknAgSTK1AcRigyELmuIelL/xTlFJa70DbuUfu/6gvYaddBvGVEH4Ak
CH4avYI68sUkPKzsOJnqmWxoNlBrlDaRnCRbVS6Qn5zKsmDpVzPFhVPYTOlx6lke8CYMiNaUjMT/
ooG3LxHXc5C05+AX4ec65N6vS9bAj41jcF7G8xR1R5n4ulq5uTzWPesJ9NWWZZczhNGQPkbIzmja
c++vcfEajGMwHFHIrXeo/vXRgkq4bVXiduDu4cUfshP8wiFF4NgF7gVHYP7wMqDG/4kLHhWdzLM5
O5iq4/kMvZQ1VnfvDUUr0OlEpk2V7thGnpJ5C+wVK9X5msu+mgZLw+9zSYMnwMpn22zlEun/odMU
KEG8BTHSqabzj9pURSazawVwWOmz9YjMAMW+MK+PHMlGYdhqxeOd7jqijAiJdmByc3ggbh1aijSo
Sje+HVlP/8Q8lkj1V1WjOmChGVtdvmAw2/Wca/5KTpn4mPhtKyKGQu/srKdBv68SqM/HF+zDqdiH
STArj4b/L8hTcTRu9kmsJpjzgJTXo5ItiGepD1l6qam1s39u30vzfaGZAPKOg3niBiR0vN/5ZkYk
77AzQ0Cx63NU/y1nDO+/Xkx+4eMFO/nbiU1BLy66kM1fbdOfANWFlSPkUqp6K57pCqtQOcsBqiPp
ZQVRf/+r4XnHmweEMzGbQA9zxLt6KLhYsEmXET7qx1MK9N9TIbYACj9JVpMCLGwNAnfj0o85ExFm
cHFLKULuBPR9Nrb3eeHIOngtYuCRt7brRva/5pAJ1q+vuaPqp/x1c9RiT0yWkUP9zfVgjTFJqOky
QAyB+XClLESxUBDWUdD6vok2WUvvWetYNp6KZnK097+Lzx2vodWHDLsYzkd8IQKoR7FOp3HPO6Bl
/4Jc+/APWFE5XQ9i7idK8XKGNHgY1UcRH3ztkDocf1DlNIlcVBZCeRQqNMryLxKgKAksV080OcQR
2ppAAWYwmrrEZWX4NmC8gzOCPk/P3/160K8lUSQr054KCUp8WC+y2ouFzU2J51zO3gMNi2PqWGXt
rQwPOrqMr9Co36ujNcVuYahLtWZE6aO6uP/tjHiF/moJhdL6F7oM00HTnqIgL7J+U3airEX3ooej
pUlaJ+QBY2lvtd7BUf+bIe41zz5FPlby0e5kGYrvFSN4t8mIvnyL80Alhz9qq5Tt77CJWD/duRlx
fC6M06JPaxWWSx6tBLlyGArMAnN6P03cUJYdSp0iC+6G2bl6PcVspjJlXc8ZeEjBc6H+704oVhCE
G0xQObHPpMkv9fVPkT03/PnOHUwatRQNyrcPRT48+ivU/UOBOXC7nlO9K1SLxR3AgpBGExz4qqYN
qqZzV92uhi4CDNEnk2aE4uKTR7gCSd66Hq169subqncPoDrTVL15zJuigeC11joXY3G1nAqShaV9
hmGcJX/sH/Fk86M7dGUmd4f1bUXeAsmZnMuxQfL5tfTKFDpxrY2pPua/b3nbQvQjzmzGbb2ujpIW
FxrLH3625+sHkdVrPHSSln9eEpIGbkueNKXIF8T4SzdzHcAtozDhGw91HlWr+z4UECDhZTCAxwwr
o7Ei2tpqCs6DxDZmPWzSm+KIpOeAPIc1bFJW95/Q7vvesJzmb3Zwu5ZVWWJlCebZPTik/aRTEwCw
pj7Y8OcDZ/u72xfguxZvqfoZbWLQ4zz/zLVIGuXKLQuUlLWbeAPFATlT+9IgxTv3FHYE0eAZL4YF
7rRCfN5Zn0STBxTFxeEcLbsCnsTWnxiVRSZ5ZgJU041Ez7MG84QIepyA+6jz8tg2YTdFL/TL6rjA
oSSGd20/QDVya3UcT8AaT0Qx3h25GIR53fdGNZU4DonvarOJSVeW1nc1kpOnj2dPZlAX0i4n2PR5
qh+A/y5+9zBQ6g5pHtBXISl5LPLVDoGUpXeBplyX4kK6BLHBwETuiS0Xk7e1szm7Ci18tV1pmL5C
Gc/Cci4UuUUUf78UAmGFmPbV1d+pHDTP5rHfFL5aPeu+sdGAqXRkc1NkyDi6wX3G/m2SRsuiRCXI
vCGLVXy9hQnLpIkQxgdTKLuv7Jx6ORfqlXNzU3kiICIFFJSMKU9y/9rinI8odK6RuUSVMxbAQArB
vqeAnXBeDmHUANBpbbNUWR34Rad0lFif/ie1o/Fn3akLRY5jdG33dNl/P1bnoXKorFbALKxYrLZj
ChlMJ4IMNWSfmAAvVlpIISBG/GUa4IuuAW9gB1uLtJjO0KJX/Yo5ZsrBUSiwklu/Q0KC5Ht+QdoH
GEL0IwYNlESSwC8DdNuUlWscGgg6sy9OCNrrhjAIbooingdTO0iUP5BXUEbB6Ys9RvFPsIk6RMtL
r6iqm767nIiEXzpQKhHpLYU9ilW+IfYmnXLbizCUUpvYcA+YW+IfQlX8NpBETkV50xAPXy6TfThM
n5GrLvXdekz/9gCpN8tUoOoQIGgHnS6TNcxGBoWoCJo8fcQHjTKIQlV4DbKux9MtKrI2rj0jWLyO
gUX++kvzHTwPdRR3Y79Xzy6Akt9cSIDXgZ8clkW+IcYyODel/H8ax0miYQkUa2MJVmI/wW0HZd+Z
IJCCPGCogYXaV1/qCMn+wIKvs+iONdDC6ax54jNBOA/embbznwitbKn+pZ9dehTuj+hmyG/AY9Tw
mfWL+q8vYez7MfR/jwA+9ZCBGXmmQwvdrppaNl6BIhkRRSUlRs+J/wvS6IcPghB60CkD+IQjoZpg
1+BwAejsfD3sDe+Etiec31X9bpH+nUrNLaOYxdlNcxOYO4e+7I2hoEw4kLEpjMw03WybzhbhgTAT
KdcdU2qlC1Kq7pb/MSDrk0PHpCOM3uohAiAJVn+zCg3ARvHQHfcDTTcX+fRe0FXs+NTGgAFaKFie
oydF1E+ZG4w3oTeVb+cchDhYNHVfVG1zJ+MwRV4FFnzWN1+v3K6OszRiYWOQJZwGd/DI4K15KLxX
5QkD5v/fyl7nSPuvrJ0/NzgEyYXq6RVxDdDF+cJvGHW22KDzqtNXLJpeaZoQ/aCUw7/eDo/kStbR
urPCxUJk/+Sa9mrEpLi/O4pF62wvBz+sAz1tpRbSrcJgNdbEc2i4eotkEsix4VVwzZf2624o6ZNM
e0cOqxobUphho4dSQyX17X738THbXMhvUIGqxTGdlP8wWb7rsOGLK5lPH/mUaDA4BzwW+JTHLjUU
PsiouZmpEdrVeN7SuusTeUAGM+32Mm5JjN8GGrMICSih0vAs+qbabmreVy+YRXRmgRlAmrPIM6LR
W4VC2HirZud33dOOP6Sig2SMdzm25j3G3x70MRBl3LzL13FMNL1JAEhIhwcqFuJurvTXbC+fmMUb
C7ZpKESyZ+Fj2C6deSVxKvTN+32Tk+MXsovoaVmIhCkWhS4ieRNmcwPyH2YKAiv5nqZKjLQvFNA5
rJDKtfjpz1OXVRWJOyMU9Yl6XMfMqvFreIdSyXtwvkQa6v7PDP6r29u78IGddDKFrt6b0RxyMPP8
11ooxNNekHx9WzCx0u0lSr8kgqnzmcrLg/6ArdC8R4hWwEv9x2o0Qu77ZPPA+msvkklZrnYC4U+1
dvOn9aeyLZt8u8IUtKa+4+19fTcvNOJ/dBeaqj4dadxZMJuI2eTg4RqgtOE//L2Cd9kMZAnPmDbG
R93w3A9qugJx/Hz48vzFTT5GfGOgFYowUXQdSfAAiyiLLL4kZKmgacBjsizAqPwd014IdZXVpahu
rrcJyMdhcWgTvCVxIf3VR5iTvNnNjyTrJbH357/sr2A87G9Z6+W21DPe9dmyKJlY5LV0d/SYr9xN
CrnbqwseFleI4qkU0Ka8IDaCDg3I96kihAb26o7XN0PlRcSi1AWGIqzOyXL5x8i6wkH8BtEJN0Fn
EThAR4hgMav1HHzljzwNq+10buER2cQX+RYU6qGN7gMXcFcmivE8kZFSuVhdV70jGDQAUARW1VNl
JjJEKInhAfc/bM6qIhMOeCmf/9UGbUsWKKiFSXCK/BPBRuh8js1m9PQ8HVAOiJg5p9ZIJbxXOtVg
ljf3vNMw2hsMRldTsoQ4/ltmZOJGGm6eUzPYhNZbfojMEinzN2NTGs4agBpuK4r/Ddsj7JVpqT3p
We3lmnYAxqtI8R5M0BVC6hjapO4Oek49+elGdCf0LKcW9sO+DJOJu+61GzJUvqLVL6j9+xTpjAmL
dy1eplaNtTEWXACPz4BbFkGG+B7UYm/GEpewvUfTYcPCPvyfFDhVmfJ1eo4upvBP2n+W7e6Gd0ef
Zu30IHu+2HqqWbJEMdQBWy00XQb0Z+v7qwsosBP4eACS4AMUKLyx56ZSmyJTkxHVOrt2SR3HLSHy
U/BTbRkaQS5BI6B3aJOn8VsMIilHX8f6HtwUAYpx/BNMkyFcVYvRUxBanQk6Pn+OMfhpQYnLSIz5
wm++11UOrha/w1M4goyuDJsYUCBY5tREKpxsdFRutYsKxddXU++tMeglCFMCiVVXmtzt1XMoXNEO
CVaKRNk7iCcW/n5lTxd3OH6Hnu170IzeGEweTidJodaRARIi2+YAnagxtqiSroVhyF0d11niXs1u
5ZkRnaG7f9eGQWv21IHD9qQTZBz9Pa7WRNcK3+ou7mgm/F21HewfzqS4+kngbgrLTz3ltyxQpv8Y
eZ8iQKnu2wF9+7JHeuQxiG+cPUt7KawiVoCt1JhnuuSJCWe8haXhw+QH92Ad9JDZSc9trR+GLULZ
BpsRlyDWWGpKfbtrV2czNLZILfvPzgkYQzYz08yf2IsBY/9Amf626rzUYxjG25CqYnaLlYHevCzT
A5yc+bq8iUQ0K/jEWXc/L6XZvIOO5/N+OKxMY+RU05eM7NtpzHhg2cKf6pWh62/UoYUC0tcer+Gc
wdQpoFl01G3agV+79Q1wmmtIuTeol4GBivLN5ghhG/By3SowslqwPKDtSey6saPTKqrMOFa5JqUz
8CUA9K60faABUL3x/hcEiGFbiYMGrs1/5YrBegxs22bBwIvQAnI5J384I5tpMrGjXluMfEQLvHwf
TVPA/t0DEucfM+i6oqnlDG0t4cz+zCdnHJCjFJ1LhANXZ0z5TIQofCwUBgR91KTCezhkSRU6e8++
sshfJBgL5zCWFZG/JVeAZh1pFRzrFYZGUXQSVAMooH/B9Lrx+LV0yLz1/Dgeo+m3hKgPIQxDSwXt
CTWtoC51P6ZlsgZr44M1SOL30YxaXTZVcS0Xc7FZXgQNyT0zzT7K9Ueu8KCtGIwcNXrUzyU17poy
zZSzPBS7eB5Im6eMubgeGIhmLaM5shVEI0eywvyYfSvIpD1G6fmT9aTZwwnkX0HocNMHRyrhjmCr
NjDc8+3xhzeAaBD89EsdPDjQ1hCCxugRLnfPFVOe/hZXTmtFEwBu+nDeiT0e2GbOPcBPIJojS+xz
O8tLXRLH99t7TdyMQINEhr3ZuAtl8yNEZzSK7QN9zXaJC9nDx0xg1TsWWvDg7ej2OA0/KT5EXoWU
R+ifmN/sdPuj62XmYP7xs5Srra7YHCh9FHLW/vnIGj+aIrBd8O1UE26b5Q9xRqYYuAm5N6cir7mT
1qjKG8+KvGqj4Ty8PKadAoC0hrULKnpQzyeecng4i7UnRO3IZGMLBLMEGcQb8NsozMkGErdNWDKn
nWLM4NNKEXBxtbkAsm5n53buEaJGY/mtATpsKpt2EARUjtaxljxx7vE4Udm4sNHmHhdXKg47ZAGQ
VX1lvTU3l6pf2gHUkE57SK9FqXxgc1pUdkDfEcFGYO6PjFTMmZaWhs+tREUF/dbcQcg7VN2Dvb5A
M7YraMAxsAEd+rsIcJr4Q0z+hQ3Xqe9Vt2DXsmCwTuLo1wBkxZJJ+vALeudsCUCPgVDBduYMT6aP
Yvq/vF8mps9o60OeGyV72Q7OzE6q60mZ8qmsNFUQlTd0QKsRejQvdR3fVDvWZ34J60jIEATEivKJ
yt2ZLHCWlYytkRilwpRSx3s3RDXwAX8dO0r8xRNNgKx7PUG1d2hqaBCxos8BBvlA56EPZZ0OHZYo
ewiAZ1AwwUuIkgmURWA3Kf7E58yVBJvLWeyhLtDQg/b28TYe3tT3gxAcQTZDW3s8nvFwtSWjCssL
w4H0g2tejODEU0vfwc7jyJkQ7PFkD+oXVWi6/XChWwxLqjkbWP+R9dkHdy3E659gBPmN0RILAHtH
igRxZUcAYdlnknLSXuMoSnHFMu0NrrM/Zo3rtsAcQQB0Dk0na4o0WUpoCVbm+lsm7UFLbPWIGSxa
gl5cc+Tlc1+aSGu5+YEGplM2xOYWa5hn7zS4huxORpYujEPMDUMKYGwfwxeJiOET7LY7lxc/8vz1
i0qD+Z1gpBEY7+mY/htCc3FX9kkkTndd/4yq+d2h8OzPtBSHIGL1clpxKhkN4ZPOEG7SnPVJpTa1
TgR/GqrupBpSt2ewozu7eMh522ldmWSf+YABEQHFxfeUQWsnRr1q6Rs4fKGcyehyYTuwQ5Almqnp
4vqQHDuRQoCaMoc7OMugeDe2n6KO+QAru0+ePxYWjQB7bWPgJpn4dbUNwwFANINTItvAjzEq7ZGw
tYp/hyvnyL/Sv79xh5Qc+miB7VmBTKvCufEAbGa1gcs6VJH9sA7yFkV5U6qbZVC2iMpybmO42Ri3
adKnreNKM2HOtFRXAInuQpf2YOxG6rMOoEGutp51Rt5qfpJJd9OF1lWA34536kaj+pyy89faGB++
phXBqzVPyhujbfsnWJmMBsCp8u9a5v/ugQ0WtWzDaJS3qkVe5jCN6KXFLDBQOvX9ETwrYFP2O/x6
f9Sw7XWtSGeOYzK9t7xnECyO9KAwo3Znl/nqXh0OAXHyfQou4WT62/52UVnfT3WQ6B9Zz5CVXcAc
4iloLdzM5tCviQSGgoPY+9Who74mI7Qhsz+hnYElmM1R9b0XGvNT1S67bZn2991rqSAkLT6Nsy/V
E3AEnh5n6JZaRjzp/Kr1AEf2p2Lf1IIztdo2EtaDWGPUsDvOtkh7eY1B57oJ3BGFdXS7pjwj3Nbp
KdpbPap2RqITbTrgz0PLR/6l2I96C1KxPzgLDc4HpwLGtBnAort5QMkiS8Q11XDULyGrOMIVcHmj
5oZLA+8WwntDrE4V9OVonJLByDHHn3gEDjNMgYdwNJrH+9Xktn2NyKr4Ts1E7uhL/qvtt/r6ks+7
Uy2XRHcCfouDcXBCth5wazFgj68Cq6SAmeUXJ2Mv+ybHL/0PTnx57AReoyz+qTAreLM2thgqyug8
kPtSJ5WlyCdW5bSu3+0geYS5oF1XSD0+broijXrqQbrYJoEORm1H+kECqCqUhmX6SAWk+st2O8Qz
VkIz0mEtgn+9eAA5MjBIeIw6qky1jQB03RZewkmeMJR2noIJXP7nF+xqe/Rvea9HXwmm8PvftFbk
7k/AFdk54wGgE74fQb9WCureQVo42xKQA5i1ajGnekTmSuM9ivIQpyJ3AtrkXbKFh+EH6p5nYEUO
3mvuItvEeRlonxvpsxRJvZ+9/xZenGPgr6ubLKzAqY9kEw7W7c+nEGNlgsVztv9u+zOEbxeldZCW
9aVGJLgnhF8cAE8gUd7/I0xxpBAHOiQ0q8V1j994qwS8wfFFOHOS+bnB1EhKB07SnleL0+tLHpZd
xDEb0arRtVv7OslBt0+cqqoqvEWjoU2VxS4H+wpjmBhPUan/V6egxWaScyZx7GV1Ng/3AZHMYTV1
syTyup/bt/dxzLrjZMTk59AoJgs9I9eTyg9LCBuOpjRIhg5/Y7DrQhrYVMDLIxz1AuZBnQuP2fnh
Do8dQreOt/cRwAs9JFz1C7tX2COquMiM++KsAXWyWgcH9SmcF2vzxMi22mM98GTLQI4cxw6zNbmm
Gbu1bVywg/VGPGBpNF4JKA3HNyhPd+KO8kvk91vo/+Yzs/IzayHnvqJ7OZkDbpSq0U/n70wfPRfb
l3oDlo7gvRNP0i6Y1AiKh6ufWMlMzlbddMbkOXN0rB88M0n9fywXu+Fc00+nAV2CPoOSv2ErXXc2
9j1z92r4CDw5W+KSEojPVSpG67bY4ngOx1bN/Jw4P38jRLUN7wg/xAkI4YZwZeJ+DIn/Y332mFSV
HN44twuyIrp2IkW0kB13kLJOnK91AVy2BFMBNV937rolkgdTwVovgTrwC4J85fB+ZqjL1T6YqU4s
wRCjHyFoxTc/ADJhb0/xnxbac0ODPHxipwnYoanBFS/mrqCUz0u0ixYwfURx/SWWNbNHXWu5s2CV
CntksgMVmOL4xeHXEp5B5JBAMAzfQ3MNq+1/LFpa3pmnG6/RuJOWqn1j5yu3q8PW1QhW9px7DxrU
orto0fNljvNblun0TtTrSfREb/wOHb7VT4AuOE2R41QVYTSOvF5V1MCRsIYQ3f5qbYpgD3MvuQkm
ise5hMRw0VcBUEash+QHRKpcpmZ7aL4CAE2dfKKLSU44bI2S8fsPbw2/0MdAZI1aZeTI/Av9uCkm
cNgs6udWR1O5VEaS/DwMlfDiCllGAKFeksvg67nLvabwvKxr3V+og3otwIzmXpADQx700UATPGmT
vU3vOQdMoDTi3Xr1P0CsOZD5nwJok8V+Oy+m07aLxnR7Ii5nJjHLbI6dsnNs7mHskz+E9XCLfOPK
/oyfc0I29IFGV0GOXj5EKKqffx7RFgIF7p087FcoEmXTGmfSmuVIt5QePEXni+4SjJZEppWDNXgM
b9dJ4dniUoOBIzadnty+mrNla0Bjzk8Kp1COzKA3QH0iEhJ7CKfCFBrkkRuNbmrAJq2+c238EAYL
iu07GSNGolvm+BiVWd1JMDmaV6QEJTaOivKKYYqLBNFhIWN3ywnUFC8p0SbgJUugB5hj6C7kWz7+
nVFNZEVyq8CVlqDjD0VHzgDr4GwJxqoxmbDYRAK15WICXrx1sLRkitCLkGNYR+3tWFbRSvaJMalY
BVQi6J5ACUkVoFJpqsY2ojYabFjeqXwM8GXacjoHtWJpH8W6b1T5t5C5cxl4Ia0kspKbkRbm+vAU
CB1gyvvg/T5JPnmLpkbzTzbGMxOVaZbChd7lirBImzY4ToQ/7n5+naVfME4GZFuHnWHgJ8VB4kJX
RAzrIicwcY6hdUONO89uKQU05Q55URVFY2ynHXamNdHGTJEY+YmWua3eTSftbqXX8dxWzPGCHyss
7GzLch5MNjd2Iq46jUN/VRhHILpNLMin5Rkie7HHiubVCgwjTJ9BLAh+oRnP2picgGeB9gBn+0ES
0kFU/yIqg4yIWqLAtyzor0rpLikE9AgkgZUPL0Be1gpzUPGwkKYkDrwGPKpm8HB0NQNpPeAO8NxZ
j/r5TMX0bOzN8RrdAVvDYQ4X8UvRTB1yfsDB7LVC5G81gVhKHCCUNqn+C4uFBSzfEaHGWBlNc8bL
KZM+EZxIG2pH7oFC3K8qXPIVV0uHXA4XQeQ5wT/gtR6RI5k+Wzxy8/GZVhaNFiN6udM/gWmpRu+a
AV+EMvbr4Dhaveau28ZRdq1WxBTTK++lQEucoNXLvBp2jmtMUmsOF1ft8pmQyEe3PIi0sFqchy5D
ROWyfdxYNCk5OvS9qbgffnCHGU/tcIn1bZHP1ydxwsg4PTQYrrG9+q66IP6xVhDn3dWl2tEorWDZ
NOi/Hcd77lv5kjzT818Eooa2Eq/7XwFLa/N/PH7l3JAwVp7743gclYEBbZuijmHTN6D03yoE9jV2
XAiNX7D35xG5buaXa00fHwjHaVvooQr6VxJSYSIRZ9tRc748hilTUUkMlF9aqoCbvesh6opWwpLf
vkK5ByCMagkDVL08TrBZKvgrUDp9ph4Q4BUR5Yi8hRGYVMr9wLxLwmAhJfEre05HCCYJxBxomyt/
Zy8JhVzxE/wQiDnY+pJspoh9soxm3AqdERzYTiz8peAxg3bfrE8Mxy3zMvAbhlzOZuRgtVI24WO+
wmedy4BphpFJnJLz9i10TJfHmfqEXchMlWAxErRMxVCWlTfj1hZrBqlr06M0KvIDd/wfWPIkfc9g
Rlb4fYTp6RVrDyZYeFUPd2IPfM+vv9C5rhuAaqOAnhjemwbYWhC7njJX/HnlMgw55FURcacqwdba
LJBIDOD8fbA3eO/FT1fXC7/BCGjCu/vQ3D6rYZjwYstJ3fZ3gEBctD194yBd92TsLUIWB363e8Q9
L1e+utl7Doq53gDacab3j5rd9uVyDFYdu1XIZnPIwG9RZeFm4z5Uhafa98j24wYxKdANKl2skaY/
ZfiXyWI3fs+Y6tzSOaSCYbatYU0mP7F8qrY4OzBahef2/qaitCZuBK2AwPjIr35o0Watwt1kZj04
St7tXlgaqo3wZm5iPClFNO7YD2W5jKIsU/iojUMEBvE0+jsku65PYVk3iO6t7/O7NXXKNWBIRGnj
MuwYiKec5I5EfV+pvDezoPFMX0TfUTxTj2v37RjTaWNqa3HRJ+0z1KVZM3yF/B+VJx13e7R9csMG
bNlc0dAiILk0u9+LICuaf+uZjYCiAKZI1HLvJFPyE7Qdev69WKEfb3ZqWrFfl0GtK2suy59x8fnK
bJqgaTLTyCFbArmuVi3scVsmynubVvuwO9j8ii0oZ0EiNCeq165w1XqnL9ANYZs2eFLzxPZ5Zmpu
FXRSLQYkCOd0fJMfIrHQCveN7MU2kcslD0V124n8ybFOKwWo2xMq/m+rd+ps45f7SohgP9zZT1Lf
Eg82Sh4JIdmwn6qvV5Ic7yCuryvNZybkwqBX0YIf2Nh0IL1FVIe0GJ4mOfKZHPaAwSUzMguuRFeZ
gvYmL/3L8Ne9YNv1wiWPDrCn+4ZBjcec2Wa3igC6qV/AxQ4abRh8+cqIgQaaLgLMhoKaArJ0Y9TA
TY6rubaAkxplZkG+s9V/FzLYYNTbOG+7pSM/ICaZ6r+6YONG1o/iSDBM5ImxUUjw1+vV9QF7j7N4
akqlZ9NC37lZ3Ki9oIuPKy6qdIq1icRinRzb16oeIc/K4kF09MwyRfq1i3wfNTG4E7lcT+WeS5rc
mPEvk/CVt5hnktvkBREtUnAHdm4TMxby0I9HqC8MdIcZola0c1Qh6OAyYm4T8rQleNhpycWzfKZ3
V+39HS7AautjhVf8ExrqEH/SXOaAPWlCdGdBwPYTyu8I8QP+WNkim7s4IAZpRuHvZkq1fz4k7uKq
o+5bUBVHOW8NGhLCMKo5lN4EUwin5HnjC/nujIyzEC71GVKV9uwlyYS8CA5igaK4j3QIWYPVdRSS
U1Qz1MXl6P1y7aTRpWR39JbAKDZOkxhNFGQxwVCD/z0qbnCYauir801/EJMtnYi3o89Xzqjk9qeh
KMMNQyU412Pfspzxa10p3ryCCQd/r4zuUE7ibU46ydJjcmvcZaDBgU0+j+ISOeSC5oaoxsbNDbzH
aaC6CzPu9PSC3yfSsnednSVlHjHP476Po1BrJCPah39tR/TqvanF61Ushw/t1fLjY2MmiWPbgvkB
Pv9L31nqogqOg5fc9y0lbzYYoqVmUEisaht+FjpCsvhZ3CXix8z4zRD/1iMCOueE0/2h/eqsqeER
189PBahhm49tz50kViLQLLLj0tp+asHEaNMET8V0gWXBAizRtYXm7EdA3E58XtqJ9ahNaTO3Envm
L6t1qnToUTaj4Kz4vOM283SvvYjpQH96BP5qDHoaBygUSMENgH7q0OltV0fv4GEtKkY3yj9HPk37
nz2iS9ONpjBzkew9PtweA1ROhZ4+V2bG0c4IreHrI4BHgr1kFNGAoAmC9eJiGOhvcImQrvBPHd24
UAe3X30qohp75wDoQ3BUKet8h2mpXw9VbZ8yQL1yu9yoS8uaWEWDejtDabpbIGSobeJCbrtjTRAM
uLgDpBy/EJYvIbur5qsWPPibPQtYLYmv75ze0CWu10dvrc8scCeVqJ2gDQ/RTFiq3/nW8fSLcvJx
0/7iU6ozrpWF/jbXXzbkSf6KkzjbuCmaxfK01HzP11WuC9nAmTxjBY82wdtsK5JBRghHPZlLUt+c
AHzPmVwL4f1SGYa6SIePjmnxpThMVz86gdjzzQQYIjhdB5ZxAyB8TTGIfEkAwqV1ybty1dBnOhoI
lkrG11/g7CApYL5Jb7utbSH74GLvMh+MGt9z38UyXWEZP4TzwJTZahGe0oS5x9JM8xUnz48K10M3
MSB9Ir8MNrJ7+uB1vn9D+5c8XiQ+SjrBROeEG69JsV5AXMC6SC6XS0PYv2ixd+msD0F9eDvF0Cu0
aMZ5KAfc+dU3OgR2AufkntPpC/q1FtFuoL/9vXvuLB9K2DwD5qfEQJppB1LZM0bQZJD/6tELXpPd
oHZnUS5wU+DJOk9z6a+wSJ3CCiLAmaY3v5Kyr2D09ctcA1L83XVpJ9cXQUpMK0wAVrf+D2SUnZzA
7KdVkAys6jSBlqZjFFK4dTjFSc6/dDUsTXnu8FcOLfYgNCCJAXUhKm5JSrl0dlgYGYvmZs/4mCMJ
Ai9D1YIZ3tpKMI3LFXsZ38bWaMiSiLBKS20kSdCUQEquYERsF9blTYyY1sloi6dM26WoVyo1JT6H
2fjnRbAytVh+1g+/UvDFQG3cVkcVoXIpvHfWYXsetOHZR4btqKOunjP4iwN35UA79mmM2+y9uWpR
Ky9ZhXZtaCAWZB/Kiv9ws3tMNpX+bYYxTmtzi8BTuX86NpE10O2y8ddpyO5h/GK4+fLukqqElM0m
DbCQJp1GpoaJr3f+ezKWSkh65uypmAKtIyMXQpGSk0xB/s7wIivrYP92h+K/rOAtb7KFdYfxNNjo
q7+ZS8g+5Z0i28lrReuXf0wtxeRzTWgG6mBzwyK4a+PHHNRsIrQuiTDV1TGDdbRtWeKKYk9x96Ph
03jwoxKR3TJovGvL4WhmrdavLVXfBBxwh8FEd0ZxukttH3NIPyuV0vawU12sl72HZS85P+udj4xZ
zKY0mdCnFb8ngBq83NLoVoGOiutoZpjINsAXAeLyTHb6cegO5z+iTPy+AOTxIsThvJgJINyYrDD+
mXm3cFiaoJo9vfbHsSFGbtxRZ+PjL6ssAB7QXqUMuXpMUitNDlA0eH/YWYZCwx6zCPPJG4tqFkb1
AHyjqFv2t4SLASxsN6rJzXr/YYiMfVPo1vBU+zbMROGCATMd6RVgp4p0O23oYHcPBH2pleW3QFyJ
64cJgI+PlSd9OLPVrFSBaRwZJClM092EzvCAltDa7TpkOT9ZlKKIdYoVIbys2bTLHBy2TiU3gP7J
BbMCT6XMHwmjLpe1MRkKiLlTb2emgUG7zfrpZLrq7fYwAyD+/7gK3+tL4ljQMO3inRIotrAzTDDs
GwE/WneJlw7z61k6gQhqhnB9Rnp6kIhgrpoJYpTdv7xFYXE/4dUmsJ5tVGuPufFxNWM5rZoEB3N6
yoZ2cD6+TIXglprQ7OcH50wQmKHI5UbKnKxGijkUwj8uj0vAdoXU4BfYC7YclXeuO7bkyE5fzilw
tjvlquTtoFz0bIfBjFkRRYDekPKy8kfwLIO1l0/1rnaqXdBqoNR8Rb+GjCrxv+lO0CLIhcLbQvfh
p6CJ87j5dJa4RKBGn6sQ1gJQTeyv6bF6Q1OgoGMzdcUDzy5mrvWnnTifoo6iHkkKC5wYmvA8zdHF
k+yU5wsmUZIEUl4wqxlQrrtPYK0DeTlpgJUcF7JSlJMo6+Vj6C3j8frkyODpUyE+rRgsGKJflZqD
xMRhgNzE7S1fahRXt1OE/vD5jCgZUnFNlXkROOthvt+mXi8dna3q3LFn8wWmt0T83F6SADmEanDV
yNZ+r79OntGFZmFM/0BdHG9C6056oqGFZLSsn0LEcBZdljFxA4QPUCt9R1oqSuBRANIlbmynd7Lu
bWMFa+ECfhSWr7veQv1H1LmxOCLzI+oW001XkCXqm7I3xWpYX2sEb3EjQqXF2ADKeJrpNR88JTJV
9l9IQrNbDnA8ksGca0E/H93ozG038MfEuke2iq/lWSDqw/fu+6QfNuyaGkD2BGM7zva6WgZRLxUi
ixmkGYrRaR14dnNu4qFU49lU8x4R2JOeiRPGXdxjmBbVNQ+jfPBCAYdoe2rYvr7BnxGyTVw4bFRy
Zx4n9JfxDcUg5jhVveJKd1srPgS4mOoAiEdKnBD5ww5ckQoFcN6x7Iezju2jelFAvYuBAFPUgH5S
c95RSnfw3SIWn4z+6SvjIXSM7O2p84oxvOedwZqVBXaiwb2EXSfxrorYF7dhI2icm5XdMGsLBEOC
d5qqHDGQeZxG/myoz0jLN0NQyKJyKU74xSAVPe+XNlUPnZszPhcBOV/8EAn6BHXFFPzDdC6lzYIT
IO7eDKNju77ezrbHQBfviOJ2/ly5O+3vfnueyQCZ05EkmHGr/ND/YUnlTiUWsewq7QelkzrKfWbP
5xzDCH35M8FYbesbdV8N43jIdpQKqYl+dBDXrp2IcY5TqyaTS0V0Z7INpQpJ3n7EunGZ05nqeECn
DqNVcrDqOqJTWI46EPtaA1IJcGlLV/ASOdVg0+BlxZfsLyLkm8uYc5IaGS3quqm69wxGsGN5VfcW
lFl+gTHONQ5wfq+9ikch2Tvx3ubJ6SgdyteuPAobuI98wiP5/RmBL7xZ1qvKj8xvO+kerDczanM7
9jTtuEWY3rSLHhRx6wI8jF+IUAv3PAy7NQ9vGaMvxljTdStHYchNl+H/PyRs4fVrZgDjWvg0tOQx
QRDLLicXMQhunvVAZ5HFGHM978THoam/iHNugqqUgCEU4slQq7fD2vFGl+RY6/9fPMgoPmYptasz
eyrldYYu88R5PtLfKFG9Fm1JxYJATkdr/tfa8q6gvzFj5Q6ksU5+vlnkO20/p22fjhP+A3aEXXoD
TngxAlktL8vMYr4rdSGBo2IYEuwuXfesdbg/bRV91kht9rmSgwjYobuhoxZY0If2bHimnA/alRw8
vewfgu2L38bT5O5VubSvvamF9URTjPT1z65fFXZ/DHipqud0et7epqR5jG7lr8NPgzNN2DQJQ2R8
ExL25JNUM97Eqm6xTj9LdcIHOdeIEvs7j5IZPLJ52I9Fy3t6uurazHedB5VpPwy9NW2WPeUmpf+L
SvER0qRj6C1lqbWPjLz5xafsf8CTgTflqIfX8Q0Oce7HysZVpD0sgKh37Ev9ZqkBvPHcgf61+tbt
wtddNfeVhVj9XNFulAgYCmB3dJ4N/6LUB5QVSVJZ/ENSp7RICBUmhMxIEeZmEmy77aUOqOhIA5bE
XhKxYIQmuC+6Nf306AeQ6lgQ+nEEBOiNf/NVl4uIPZv4IYgRoh2HhNUL48E+AlAwG9cQTdOy9zRu
tAzOKJWVPlU4mnbi0ViQk9WcRph+2LQEBvHY0llvLGoq7FbKbM3l7BxzxHf63pHgffTknphiJi1a
8oQLISr529FBdMmEjwVNt5eX6+VPYfKNMay6H0Rwtlo8Bj0fHUf9dd99gDedrYrtAlAId5Q3NzYF
m+jXFKvcv3Y8hxhm6Q+/QIRuXr05hg2vOFHwZ1lEzG6Gv66QzDX10YY7fUeYuU1dY00IHUPv45Jw
N/tzZ2MIHldYs+IQTpKn4YgFeQBdy9nsO2C0a65r9xqOXkLv7q0m85UIdG38NbJxrW0HvNlaR8nn
3bQvDdXXkJZO5CWatqGYxnm1DPeyoeliw/3y/yotHy8IoFzMObrPi79oUCcTjJ9EBRxLdyv77OAA
fhuww6hjIOu8MmkEH1JliZ34Q7O/bc9Lz+cMsE2hyL4gGS18gisNimGUoA3D9E82E+yMLUVCWR9I
6Z9dX+WGyp7YkuOcVx/l/7XaBXd2WM5ZsZ7dPklIzIlglRHrja7TwvRi44M6q1aDpWWJAmJgftma
vfZjzxzGBZGSFCp7IaMYAz9AcxU1IBO/QsdRv31jK0uFHcI7Zu2HjGHmpj1yrq9KtlRUe2azEeGQ
6bgsiwmgw7i4B+81N55ULoIWKs84f5Hk1fisNdrfjpL5TcmUV7Ta1EyRE84H3ikVO2bFEHKB9uaE
mZatwpsyQiBvsDphMgbxRb+lPQ/7rpljBQuZe97hPGDfSiWhmEhEACCBrujUKH/YMXGSvMTWLxk1
vQiJtQFkJIFovjWnkGpHLjVR+a2MYcWLCPPoqgvSkJqjkb6UBNLDBlm5Ug+9SXeu/pdDGMBMyTQz
FNfMxdihkSFwQ2NcC/U4Nc0xPK3Juspzi8VQ2PbRq/upaSrPfFc/6ebPoiBQYvusGyC9+wJ0z2Md
Am+oiWQ2oOx5P7e1Lx++2yyvIoU0ge3Dzu2DQLL4KvPrVFJqL33MEx4bpjw4HWijnkaNvM+VYfRY
OmTZ92/AHTmNCd0eDY3Lp30iPrK2VC+ABH6KpVCL+bmMTxpVLAVppcQJMZdYHZZaEI0gvw4nMVny
cBKaYXyjoM2Pa0XLNGBTiN5E4ZOB/D38EeFli0tn/ZsWpRUeM9+use57YTD/vhdhostvwZ9AryxS
lUcHunQGyS5gbM1nkvKO7ZIU9C5D43obj9TY+WHltWgJnRWwsYUmTng/f+uRuIZw6RrjMafkqUOl
BqzaTinWVKWb9625L1SJuJckedbaalJCM9F4frYpTLH70dKMceK3BWlIklE16ZC3yNRA3XwlnAuR
Ibn2gX05BjKuQjA/jd3PB9ry7yyW4dupG4b39JEN0AaMoTVqc/85gUmxpTW+Wsav7c3M1Vx3+Iea
32LACkQQ5DdZGdMFbsqH3cThcPEI3LAGJ9boBNdUCpbym7mCWO8rJWZzigZRWQtf/FTZ0Y1tTHQQ
0rTwi9jLCx4+Xon20jhRgoDBucv9hFTlcJhq8g/+CKZs0oT/hiuE3Pl3DK4WDI7O77KqOp0lf9hD
1URZefZdYP/8QVd+FhGiNfJaKT/xlhLe8+UuQJUMJh0RHkJyW/5MJo66peqjHDTq0oAJkMf9VeMb
tFbIy64jhaW4oK3WvdtcThOfpxWzgeaHbz4EY+01PH+uYabIzCd5Q/1Y1Dlpxue8PNG1I/2QFaQZ
hKvOrvHEC24nL/wfuqS6GQmP6oqhfr9skMMIdhEH8F529iVbbQajqTujO5WTemrQ56uqaW5WuhD7
mvSfw9Z1rUCd3DqzTO/6+7G1pE7Ipe6Ey5kip95tT9CcgbxLF2er6DVRR+dmfRP/PJDojHuO9bT0
g6mc8M3ZAXsJk6EWO5uY+VtHSS8JESpf6o4pKLxfyRo30O7rTGEcHCaGi9RYqukJnO2J+nHzQMvF
++qQoV+SgkqSwRIpHe7LMHAsSzTi4P74hKOuCXSqSnkOijZy4BjWsksrVKnn+jz/wu8XD2Ynwo+V
8EqhRuZlsj0/N+SGRChEBGKgGOl39bVLE4fAjt6hGj67d+thIAOkqlm3sbMihr6ZXw4cu9cmY96E
75qIvyqflVJF2kppCkm96t/Zu+DnugPnSgEKKsS9EGJefKZDcxG/qQo3Dx2qSTGC3q749pkBYmxG
GkxE9n6rO/q2Pv8kiRmqXutzlUjGtFJUrr5Xoy/dlxmzEpsbLpWrMMi6E48CqvHzqH6SenIvurjB
I8lA09an02VLWEI7ocSnNkpvqwtCAhAOOdl/ZWZ5mlpJDbmFV+++Mt/Lzx8nUT3BdGtir5YcEjFM
XP3qil/RzYwDnS8n1fizkz/tl3/9xYR7A4T5cvl8kUoZ7WngKuSVCvl/IDOTodF+ysDohfbLaHQ/
pbxQ1O0aR909gNR84oquehVf99lzOGoM5rRHoIH1DRj2qUJ5EmlwWH/AsvrZmum0bclwTZ6B7fJG
RbNnBve576pMbPTjkkJ9jtQlLjkcpos0n69zattjJnymJtcsPdXV/XNpynvZP2slkcmkGJ8NbzDh
oEwKcKsjnv08aoM1BIJH2zwCJm7ks7H49O4/dGDe7ff5Api0VVxp/OmNtxjNuTFwae51SG2v8ds0
pVmRaF/sRxdKxFrdwmV4/rOh3v9JNtS1H3oT3LM/sVAa4R7Xwgeb3o7opR/qn3HuUgZcFo0gjl18
KwZ3u5jE6TZj3G0ZReNPjgiDS/qpUkHcdWellwLvCGbPs8kM+T88RTo7YtjtCCrvyk48gCZvx1sU
axOBEen9HFfF0bJdZASZq0XPuG3q1cmrphv7+dwvy69ndPhnC7Bn4H/ocyUJOZL0SahFZ1ou4I9e
aB3u2EaJVHbo2Uvoa0SdplV20pijnIL6217bEYB9gJ2lYicm8zbgYa3D4FbP9vlfd/aU4P9/zP/C
6hFclPrjxA3TQ+UyfUPvOXKv6fkQlybqKoFcAerTd6+WJuuiq9N2bt86BAerUe5559dQCopMUWXq
yClO/eadFBh4HTk1JXb5YLDOvfIhZS1ckgF0oOo+EubVAB0SpVYbDCWOcA5/8v7knph+JK6J+GW8
2mLeTPsFhjpAGoWsxVAG+sm9CplRJUj6N4NxMQcXfNeuunaUkVIJ2+3WUQPy4WtC0x47j9ov7ZrD
1gotqKgJHm643gNDNpz8Ot3JFOg5Sm4xHdcBM31RuXSU1zqFRyva59+6cOgauExMOaluhP40Z0KT
Dfxa0N2SDAS+CurV+6vJQQyiNi4KE0C+TNgS9uEgTms0fhjq6bja5U1B92A9g0IF8+Xje15jtw+Z
nXqgPZNIo2/4KZF3i5BAvPpIRVi5LyFOxJtWSGLPzVqstx0N0GjggauExmPEam6LIc7tXSSZCmco
a6RKs97HgCbo1k3CRKyDcrgk2qWIQ1OlSsQEv/JqkE4qBTwJ3HxxBHgFsxp5/ypDpwyRzdSEscN0
DVCK5ngGHpdI0uf7roqc12xqmlMh/Efq0HCVEiI3oGM4DfGKYWSDc1IhZuyebPgOUuRs9mOzd9p6
ol4p8+iI2x8RMk/TVCfXqInep41c6wvZXopuYFPNTuW1jAtONkZfDt5Ts1Vg/AZ+6I88QqKpsFvc
cZBwWRMascPeMk91qShghmtGjVziwmBPFS6KLSu8aGXU+e8qA1eefE2GnrP48xoInHwuqwxd/iHl
ljRIMMlSxCoYWZECUTPcd4teI3Ib6De4S1FFoUBwv3FS9RQHrxs2XNp29UOd6X+LRojORv2KB7DR
4aEKHULqSVPc/obe1PGCxfrPGOfMWJxL7OCd2kQ7pVp5zseqUcm6ShJOOMarlI+ZJ3raJ56jELZM
FymnKS9ZLkmANrDf7lRNHd8CaIItkYw2YJ2Oy6MlKZgcY9UWHfWY71mUJQI3UY+gJohPF4NvRySW
mH5RHe7kZ5OsLCSgP8oQZ4qkTHzdgGvOjZow7FdYKsESqOOCrZR6uwOX1Rm4ByCINQetWCQrJg+X
FC3XPxy7cR01/jKxdmKXuEJTAOSmfyb55aFZ+fgYbR78bpQ/GY0uPyLVn7tsJ69NwGZFBCWzRC4u
l18yzkLPql9N9ONHPiEULfqXZJXhjVWT0UAorc3xFG2C/K2vwbwI9giwFXvRxDghPY27EBG76tM0
zIY3fLi/jA7I63g2PEp4TgEplr/hXBA+ebKSJ8wDJNiySpLxozE2E7nSvi9n/ztw3R+ixOmLDy5s
TFkD1UyUdodDCCszsVFjXJNjkxhuONW7KivD7tRie1YvSL7uIAV8xyh0H0BO0lpPodebwCJWZNU3
LlwZF7i8wYYENei43CyUpO83BkBrgiDUsapJzi37An4XvJWCgFQZKTkNpdKusj/itqDsOTYfrkYn
SVeUPAzoRRv2zCNpkCg7HcaYSNjOmXlTJovarFswu+QPuWs4EU/8O6+kTvMZbc8Dy8cC7+eBGWDz
Bz9NfiTHdv/ZGT1KlWkM+XMvXz+FVQEkRWiFCFGT9jSUBbKud3MoIDlrFGKqn0uV3XX0sq/iqxbL
5jWb/8Og+bWElgo4XyxespO2w7WU1cl9ZT+0A9wLdbQaVFLl+eC53li6hpURIL/vT4ZCfgQw1Iog
b9fdmZ1MKm9Hi8IsiZ/t8BpcI+aYkqW+2oXVrUUjlA7jOyV6432jamFPgfJ4rMN3X2qTzU97hCnH
UiKUG/wfgZOk5hiWZh2kC8MJEPNveC/7Qzt1A43OjA0JRyDR7FoKgE949JRyBZpk4+GwqCjmUbcW
HaTXzFQEJDP0nqB4FCM5Vr7SHl8TQ10iBms8i72iArL1d0HNaT4LUFrRTeubCoEMWsfE6phGZtqz
Ix5OtWUalmPJP7CSsrSaHrgxRYslqYBs9b+WB6ttHaWKWurxNq4DeTse8k6ov2wRs9eONloTJrUq
NA6DuDrVlvuBwrJUsI9rKna1uk+0Mp/QnFx6QlddHlz2hOYdKwDyvt5gZRVxhjHrrEe7Xu3Wvdjm
feoZjEtd8aUQpP4BIQwYJyOkf8Q9AKd7jidsUL9RLz+77XOOUyrRCi+skhg1r4Duc64KOdsDFQP8
gcI85TYLAKIvT11d12gefsg5XpOq7zm79+OpbmpMEj+IcqGeQ/5FZYJgZlNUwb/YKfWA892Z6X5+
IwoYS1ZLc05W0XvN0kewSRXkwPFaTjAGd6YBsHjpR4vpGHfcmEvDy7oaHuusKNLswPoq7iLSHtxz
yug7r8k5gOPteKcdKA7C4H5C+xDxa79jhgEYBAjeKiyvd4bCxzmOn4m7BFA/o+QsSrGegHf8nzin
0NGzUIVaXKIZltpSZgZgArm86/BrOSh0FpybDTOPV4O6x+u4v5u/XlcyV8lCefuaLmF1TOcx4GpH
cP7T3GoVusmAqBrc/AOhy0+EEbyVpqGyOycbgQozPzN+8Rj/Iw//WwRH3myJ18JaBhrul9b/HLI8
GbCerMOBPry8v9IMS+qWFqzDfNZVtB4HYzP9DKugZTnWT7f6NQzPIqy8LHdKsh/mJlAO3/72zEfU
cGuUd5gkM+7v7hRg7td6OkfqI0krJpMLfTpIS/+fI4H53q8xLiOiUz+Hlpuj7ahtYYafWHU9I8X7
cnXtK45Dxt4+KJzCfrnS93hBzUczbfXDj/1wDtIrRdzrA0zfZW8MEHXUPKAeeLhydaA9h0Jj2E/d
TCxjmK/YoL8Rcvuym2KCmyooPgu5xTjwzDIjexJzKFXmHHf2QkjhgveGWY+1QoeeOrzng8ibY729
IgkreJ1bfHz+iF7WTyHRD0Bqn8tONQ2GPjV95mktSmbJUtExiaOEB+9/HSR5TWH5exIIePpWASth
ptfe26Wt1BpUwSEyYkW3U31o1/PLUVV/pSfbRAFFz211YVTRqs6XUH3A7EaVQMrGkvASqPcYxboQ
pnyyPGEWiNkx+97MMToWUKJ01+uGixWSIBjyMA3aW1uA3sk7aYhPgyh6GgcL+H0OTE6ONPFqD9a4
A6r7jLKp0coTO8KRiUyd+IG2uPYjUI2PvQm2bx2RwUmnDq0qzdGsNMJeUbvpvbhi67FLlbh4fvyb
OY8kyQlId9hXQvpnvsmYKiYrYrsIng5cuIcWg+7vCA21J4X+y0Zv+4wYvAO9p3mbZllre+ODJ9tx
6lXjP93bFPGFM4/tunIaRcxwoQa0FA6JKtgyGOjWx1A2DfeZDUorAbN+yqhENur3uCYUWHVhouZa
yCHCu0Z848aJKa+WqiEDwPmqMBrON8a3V6oOyBu9qq4FER4yiBIceoLl+vvWJlie35ry7Dmwch64
ftZFH3lGm0gKPwOL9A3GNRgbROXuXMlhj70OL4blngDJPRyIWxK7hYL8YMWpdcgRlb4Uyh3W5lJ5
1GE7fuOAG4TkoJ1cMbnaHanOqd6T9KBxwAEh7GTw29b8d0zNsaKt1WGN/nJIuFHNh/ZXcxWGKzG0
cQmgsFNGrcnwbWPmE25ZVyRZ/0aqABspbfqkeODr5MTWO1JJm3ORYli8PbZg7OcFQiaY8mlgKnWU
GsE8wTMSC/EkNgkV8b9RzI6cj1+OU2GuvAsoo+6OjAQnYDDIYBrEvHiFzCISojvHNLSLrYrYNEzM
w2A5TawbAX0nflgLgHzV/Ax6DARw4PrDFfL9s4NWBtdTbofXRO1P90FhOC0p6N1sApcsJL+77eWs
YjwJUELsC+qOh7LhvjCC32CrWGem+a/WFmKaiGnDbhEN+m+B/PStqYnsCCmATByZbPsML2kQcIg2
T9AlXLLprKmET6wCEhHfdPYz/a+EH9pb8DP+Ue2cHkwYYjkJyIT0d6ITPe2gER1sHiL/muHLgEl4
QXQEwkeOxVYwM6GRcOsn3juP5xcaXkSw5/G4a0rhCPYm/T+Pkcogk/6FtDDdWLOcxnQAagCC99w5
SLPdSBHMygrRPfS+DXFTgBGHvWmS1irgJZ1ePjd3AVy+DodJ/Sj0ttS+9DCMSQKaCyIoB7LwxdAN
TZz/D3bSpKyMgB240meQfv/Q91arbeZFpHJIVasWS8yRTxxynCeuWv8ZoHgDNhd6RgfawTChhBLk
9gany6l12+K2E1yr0lWuC7NV9WPyBe8Ol1jsEM3nEbrsPEctzxQ0cGtWyoRT31B7s7qZhiRV0tyk
MrJ71+hfsVauYrhsaA1zPYU9sw4Vm7XPSfQtZUuq2nt+StQ+rtwbT6l/RhLCSB2P2kEVUkkpMzCq
21kA19O8JlMj+9Q72TpVkV6KVjC7+WCRZdG7g/fzSp5bZw1VE2uoztQqrJKk4ZIf2j1sfHdE48gP
bszXNbHZ1ioyxRI+2VY10V+IMNsOuq0B6QkMVcpjW8pQeHajZU6Eoey5+WLgJGiK5z1XxOcAfXRg
+ifG9HKog3FqL4dXXbcB46hPr7HBbjEKaSykFp1Rp0tr9v04igvv1JxUYOQRscSZKS22xNkg+9GL
A1vOgAOnG+BGryKzvOiBWyLyirW9S7rwGnFbTSCa6x7fp19aA2MybNIWimgeAjc6C2OBtXqetL5U
zbOSpjNEfdJRSN9NzYAs2xLML0NSEm+x0hvTrAEr5piP27o8TBKDXJj8tGb2UsKBH1uG1TOIRmMr
g1+1it+uw04MRWLiwys9e01ohJ5gpSvecxMULOH8c4lLBTFHRGkQ7mc5D8EAuFioPnVw07VDQz7s
AcodPiJ/uPLqzOx+NDPgI7pMMPvaM/0uOBRpeN+wdUteU8wnkpWxTlu51HeKREjROVZfknxfEGIx
jlxpUQfBS3qjCLAJodV+jpKTZOB6chHprv6yMlJPwNx8vXaN8j948+T7iZmG3s0Q08hCu8Fa2ZT4
80gbaqSD4mOXCwkyB547o19SWw3BIE8wbVWTj+xppM3qDDu+ASsCHjW76E2lAgFc2b+oECmnfn3N
deS+9xbHZvndOimIHpI+NcsZkzO0PDlOqgpmH+e1KtNX45pTdU3EM1/H+tNovBovwh0mcEl98lLF
zzmMKOSkc1JlCk7raIEpeXDbk8zuaqZ9MzjF2KRitvNZNdBV91vv1WzRHaceZVSRcT+5rO0+/hdR
ZxLFbXS8/8UoD4iNuqHV156ZnVV0B0lzaKiqhsTsKh+/P3Yzqdfi/l4Ht8b/SkxuiM0DaLN3/Aw4
S84K6G4okHnPS1a8xAmqzyIqwVGOrjnl4qTjYjZGwIJEW3i3WnYUdjq7rxmqf6sFzo7J/GpxpnXW
lACsQ3xn9XKIuBvegx1eNHDWMIOt0UZ2Ip4QW9e7Dtm+lcJZAwW0ongUm2lmS+jgPSZkVTjBXufI
XPesBqSsA7nx6HpLtSydL9HcvsN7Mp+zwFsSZBX7z6CWdSxl+DaOJDsLMVh5VPQsG27rUnGQaH1O
hscA9wHBxeJ5FXxEVOObHMdXDAFnoa1cXYoAcRifR+1YFDoEB8t6TWlIRLM4GObLQvWZiNgmAIs2
3GfljnjZjEtJ31CchP8nknCRZ+poul4x8ehxxvt0PPqgnOnAmlrV8MYQL04qMAaTysgZUNrByJS1
Po9LSs6lPRqG6aUPJzSsuWiRnUIn01ywFvSclJYM/PT6ShE86cNcodtLKNmX2InUdLcrCIzoj2kR
Fmfm1JfYZpIFRc840u5Vx3FRiavqYWMk1xgbZoG9T3NMVEdaqTeJrcQBqlS27n09T/jeDimXpXmJ
sAEJEG/1s+QahjueftvL3li9UR7SIr82fXsL78MFP1a05dEM7YyyV+gkyynXABh840aYf3qlHAUO
XzDt31rMTblzOOQeVOn2qV1iz7h3cVwMZxsstWhQ8+3s7VzMGjyycI3QX83OcCU8pwTjwHSROr1B
5HNCN4e4KVJG8qiwzZpTWE2ECRxEFSq5LlS0pvYPzMc4FxKmeWdzGaZzS7K+DYkJytCwJSlmyANh
jvjZHD/P09AIwsg6QB40Sz3eQoEf8yNLngWgqOLKQKjG8BmbWclOYdu5eMcA3dGAFN7sPlxkXb4r
mT+gxeOHEHHfYqr89CGn7cOqS/TycyDx0he98sseB/kOEjZGDb3kIdMhAQZSdFK4ecbq+2xccwpf
nSuAkgA8ntBpGc4ImCb0YPJGr0YQka1vMVCgGwIewJIFeNO7dZ+upBXdiZqPK3tKNv6b3e8soSU/
tVsLSqKt5QlYjrQ7WELR+kqUbw/K6iRke+TbRhYGuSa94jqWruuf13Ip9TT69XM2ZYZKtED9Vyaz
G/hLdlwgKBH7IoeHh/cBwr0Avl0ZtrwwPfzc+Gnin5+s+JrJdozZAGOmiVe9Jk20yjzNR3V8yrvT
OKBBbtm8328YKlu81VoQSW8OrG0EHqy7czekAzmLLBGT2y7X8ZPRWdaHxSrq9cx2DEcFF4jOrv7A
ZpBCNcbjU+EHkGUKqqcth34K7LH2kltATjlVX6vLJIvmbmLkJPMvL9Y14WBpzORjhTMOBRJbN6WI
zTSAFsPzB+/hjGjvZSqdcMz1XCsQttKRv5ewxiKEU9DxCK0pHDw62G6WvQVClJB6EBzFcOI7FhpU
V9SDKn7ZrqEuIGkoH+r0PdbY03JT6Nu51e7xq1QpgGmKep6NakMkKxfv6asZyn2dNNnjac6YqxiM
TDgAa1A8Bx1GZfAtKVe5zgVBek+joEHp/0qi7ulkh9HDJyjCFeNS9JNgeI398A5AWxyNAowdg++w
0Y8o7UcOCnL3Oft0hkELjM2G2q9ZUS0JHyDdvzbhg6PtX/XF01l5lTzYA5T7Ty7BqMBlAf6EVYyJ
pfzhGELx/qOye8CDblFz3KVz3Dv4mel5hLdBTM3va0ey2pUFcumjaNZiny93jDQ6+QCHPPXv2yI3
lXacISkYFXotEwQW3QhYNnAKTXkBGYkmt8b7mKKpK6ZcmL3qsJ9fchtmdvYJTULR2CWvqTc2iTlU
MmLFDXtJ2LHLv2qLRZhJ9EJ5Uc9h9iWVWfNkrvmoSy7fMm9cQ2O7P3XIow/vRGyPDqWYrcrMxqmF
OSUMJZV3WCIDf9B/Gnp9qyrvd2m2Wz6Tkg47IBUUpxEHbmNnP+JHghMRDpiS67LxiR+L8NqpvjIZ
RWyuAnRUEqvilILK3p1DrpNESggyln5FB0pZFmQbHFRwW+p7weNFH7GDOECsGny0ov6k/DFcKzBC
P3jMbL9BqMCfabEQHiSRtHqmctBDi/97neLaTUsyExzpGRNd1XbWUex3i6DUBQjNuHp/fxxUIcwy
1Z2VpMgh0uwsgHK/6WBY2OOYDO7XYXwSfNq98E9YKVYxrzsH7u7rIDAZYHGIYdL0vOdqB5mbmFnY
Mbz71sjaCepL6wucy4hX3v8nqqNuZO/VHuXz2c3yjtHW82j5odrGUWVlPHOYy002GiLy6f0I8THy
MGX5i8KpR5Iano4xg6hrLyktF7fzF4aVuIs0vyJ9sxFhvL0utG9lpG4d1++JFuw6Myx9Kmt338cw
/kTUV0yVplMEqgOfzUWTNiu67DqAwLtFJyV1QeLGgfUoUvwXqI9yHMGq6kr2hkXc5BByTskEFsJv
6HXkLBxRezXISVeNy5MAAIgBFSJ6zGb1I0gCk9xnl3bvufGPbaxzEzslqxYDUYvsnI/TbOKlrAf1
vLTqor/U9eV6cgLWk1h4Jdsc+44jfLyO8fJsT05b/n0WI52QoIAzLUJJ+iQxLxkkYB+D++/djKee
2S8z+Rr5IouNuW1kSf7snGaRvajnuM/gyW/dlGPbBLIkminHma5WtbhO4W0zkezk6oErw2baM6Uw
RUQVbgjDNCMGopSO7IG9RzTgk9zI6Tb1eYOcT5XMxv8Ssz4KQBMF3ryap2BYwlKi4XQ9rVUGgckG
58QoeDZhyQ0PiriDS1BKUyxv7ETGrRCUXp3qkNhZp5GIo2beGc2oKBbzjxntw8ay8an8Nl2LZG9K
LlaHncmpIKzj/vaQ9nt/kK0vBeX/cUzI2qJv1KGL/4+tD8w7mPIdNy4NZAb+oO9u8dPgvjh8yIto
VruTUgqawI4J0rTCjR+DwaJPoCyAhT5TtviIOwWOjUuCLvRQzp4h4YPygtKendS0EWYROUPwRVSW
z6hpAckaKG74pt2E+Es4yz6MoE9grUZuJqtal9nrsgJoC0bpx7CLRHA3yHKc65d+nB2wbwxXBpRr
uMpTZg0JfumRm0KmJgqVHS7nnxKH8iWxC7n4/7HNWszYmEJ6DJINJK/E76a6YitoIro2XxxDT8p7
MJVCIFNbN5tgPCnhGZqpqCdBXsiX+6x6rc/JyLNxd9Ux4R+zDuJEBaOTE2TjWUo7hBqeG+VG5Oq9
UYwpwuJd7JsdADM3UOj1oSpZcKR8AdrZD6U8f2dr6Z2RSA0l0IWowRzBOQ5MhkVWkRQ53b0zK7ih
5tQp3qyzCdQRAIn5TYefdnVUdA7hBkNMU6wXM6z5zRCmUxSFlyAB/7daYMMXsU0FEJgF0jMf51k1
iNzMqYDr6qk7zTMGoeR6osdKtL/P+AJK5QZXAQtigbDRI4xQwlGQaQN6/Y54LefW2rY8GZa3JCwu
qutJ3WadmikRrEfAUXeDeyUaIk1w1RuZfK+Fa6c+UGtpum9YPpAv3w5NsSs74rYi4pH1n6Bk2LWE
e7gLluNskaRGaXkUoi00MVwVMekY+SDT1F1kOvULY1rH0rOVdnexaBluFnIsmd23Wzo6+Y9dBIkA
05gScjGqI+6d3F6YHdXPBP8Up+k8dL534bbeVcPaJH521Diejw/HzSLXe7yVUBN3akBpqdZNW7qc
G0biwoxMMnv8U4bMZr0K78YPKst0GyacmkqdJ4a0h5gusuIDDd/F90s0ir/NGWCC+EEht/XkIFg8
wiR85cyOP/1n2aANPNRGoWvWSPPMXbrdCaLn5C0CXlywhtf/666Kmldkfpr7WRVYuMk1ctQCDRbz
5t8xrQkqeTMn+cM9ZBmOfJL6bZ030HponQzo1RmQVES+li1O39ch455lRuJOf2zY8vxg9GpKzdLx
dXoQmw+4jce8kKY8W/ZBo7f3Is053eae1GnYauSvAnVGuMpAw47AkG6n1/4t9jsl4dWLH7tmA5PP
QPAj4/6E6TvZdBcwPMYmNUJ9B3MmSPTaMtNr/NUKXLxg1oREP5P9wSibWDmvOLh4jObCgF1ohruQ
ia4Z3EbAMQg4+rd/9QXTce7ELQzvErK57Iq+eUO3dHqlYMshlHEAA318tBDC2xPA0RtTkk4eWRqv
so0R6sMSSQSplfCD8INbz03knft47xyVuF5aun4tLNV5yQ0BJxGLRoCrxp1nmdhuPxQnF0N7NwMR
TWSWdJZC0cfW7P3i1anxtqVYBrOVI6pz4Fce2SGXyfWikXTeYgcvqLXQqoED/9UCX98mjtX3oape
JnT20sn3mwnkKhMZARawiviz4cf2NJd8S3itea8DBijhk4JJv0gmy9cXmjL6Kau70vUgpe62dhvQ
S+zI9HC6D7TVKDRYVVXd7sAZOqtBA6H8x+wR7HruO5MB1e4S1nEKOp0YWcx6RpOlruAZMfgcE5DC
qsczTvegLKixZhz+RPmTtKg9L3PRMkgoNf+CDHrZdkvNGOQBNy2vbH4atixOOMrPWlLviorpkY5Z
fmWPzB1DjjI1uW+LgJkJ2rUEAaJHhLtHfmq93fHJ+7lMhBPB5flVB0m5rox95OrDsOqEeDHKbifw
Dl6mnCuxpCQCfdOALCqAoZPd1ZeDKBFkTmr+LSCJGUls6Ml4lkpg9VpCHMoabGfiUDKCWSyiT+VM
GkVoxbGZ7GJYHiK0vKu4AlCP34q+G1hgtFnfs95HjnWUBdEssQEYi58Dgtz3I8+xHUwOQbht/Ut5
oDN7J+4qdpHHUFy9T4kQMCAELRN+Zvt4QiJCpKht6Yifs9yUwQlb9G9hgZR6uKJmep0l66kEDIVW
TvDGud1w7oZXTNsboEz4dXHCrJ4LCrRbos+MgVWysQEcb8y6RPq5TyfVEgxs+muG7UqLx15pLzuF
S5FE+XQr43pUBNIY5j/GZTKrDof6yq7NoApmGrFPVgNiPSgwMcAaUe2/+j1x5xpodSXcIZClanrQ
lNscMA/SXoS02JAnIdNRoHxmnZ7tUHO6MH3MvvzM+PG/98BdVJ5o6OHiJ8l16ykxVNy7gHdmMGo6
wH1SIT9ZdUWo5oCPIoU0qOsV6RURXg0ay+cWUZNu6cZ/qFHhmuCXjDqRD4afTVU+sbM/KwZYG13d
sAajqtuH0jnBgYsis5uBYYIF1cs7x4fvi43DrSAlYrR7LtnfQLBkC0y+l4xmNh6D31eV1DM7znRS
JZjj4wbvXqwAa8k8qxAXGRw9T9y8BN0M1VPIWGjnj7zPDHVDBCoUVlw3AHyocvgctzVBxXcI/+sb
gc0mBntR1i/foHfJyolfThxjSQ/KltJdYGPG9vk0lqKKDlFatGOJGwxpJ6pW/kJGbqSIkr0WQtg+
lR6aZrCqVtmC5ogUmKHmfmXxMJaof1OnQXISUNEC8qC4ajVAWScBNalTP7flFMhxx285pEf3ault
Nqz/cM5dzC/0HROq2rjAuQGK71ZeNH3tA9s3xFNa80bN8DePho474tuJRYz+o98PqlnZiue6oNYn
RQzhCnSIx15C0vmnm4b/vQRVkX05HdpXhAEKhc/dmxLGERs5VRCcDh4HbfccsLAmYAJSoAgJ4to/
C4WkZnKXbWK295BOuJWaM816oKQDthkuFT6D5lwWUyNRZ9f9mul65yR53qoHuaAgCsLUPF7IzJWC
EPEvW8FiJqbvmD/R7Xn/VkjV4wuykVxbT79EFnblxh3fKVQA1ftiHji/UvECykOuqMPt22BGgWEh
S1I1zvQDa39az1ZCTfgYHC9apIOy5srXtrVztCLnYI7T6p3ptd613at2BCN8rwGYUCsGls/C0Kmv
TvkmfMJkaz2OYV3FFX0YNeFRb+YEpPu8MugaZvu2VZDvju1AvhfkkBxyQ3qOGIDBhYbWG5CRaccC
oWAlxVphFx1AKNORaLD7CiEYLsFOhzSjskkEoezba8QIh4nPsmX8xrO77Mb2qkL/9ot+P+tH+Fr+
N0Fld1kemMP2wEvU3+g8ROUDBwoyAyoXS38JLTKdr9gd7BUwCbQM+f+lOz8ZlRjcZFPiKkdSEebf
Hv6JZj3RJMMZh8fHBZ8HILXBA0qe0ApAtmlt8486DUxm79EwpRadQ17s4n15ax/KfZ7olkf0iqsp
f8N1ld3q0Fyj4rtmAQoBZ39uW3uCjoxLutGw69JIK7JVHoxaH6YN+xFUd2wh26U6teD2kLYKrCnN
mMFX9jY6tiwXI5EerLunqoLvboLpXS8kONkKZoPOSrQn86Lew5dYyxU3Wz/wbuTbClyps95AlJhM
CcMNIpWUR2JDEUhLhZb7KKJP6Aj0FpHV40HPmCmhcDcvw+xtSH7kEXcEKWUaS6nBeVTV8sl9p6VG
BTQCYRy/iDXLfhMbPENRipuE5lRUPwTtLXTMNO2kP2wfVJTpT1Xf7FWpPvaX7ezep7q9X6TFm5MS
33vP3PyvyaLIb1RvG5W4fLBWIKKIAZ/AvKc5WtAP3hg8o5XxRifPNUZ1o9q9IaaqTIGJwQnpR8Nk
iaXWz3RgY3HwAO0SG6OOc5ss/OdAj8wduNyFm8R36c9k5/9E7J0UEQwtQBqOvIxCsmwNPuGc6hc8
SrVJOMe/MHnWrrhgZAUaun2Fhp55UkQA6gb41pVnkzDL5m4AM4br+EiSkgQvN47H2qI6NYY8dY/Z
xxV/8j3X947ObtNIm2YpWpw+1DXtTvtsI4xZZ6Z/DxxA6+ohIyLBGp3HbSTZYQQCj90Q9Cm3hJ3L
/GmGi4NRrEtI6iTWSBhdNn4Ql/Czn9HIxli+DLFyt2ydAMpo45kwmXGzMte2t1FAwOIjldKiRsas
v26C4TMt9NgkEIATQSa4N1kgM/R3ssCZn136Z/y/EnKoYPuqNd6Nfh1K8C1ytz3/zf1gylKxnOYD
a7A07KBWSq7RfgDUWM5m6zZB+dZlsHvWgjtzegYzxO0eIrLyMVckM6W5qPyAI7KDhPTVG8ZqsDRs
8VmjRV2jwu6gX8XovqQa9LwAkB8bMcrK1jEoRpXxFLe1nS6aOV5GJ/Mn03ww+XR3Z07pymXcx8zS
8a00EeSUITsq4MbjSmVbQrUI2nG834bhlyuWxf+JkNbBfgLiU7APks1ymnUa7NP0zh1KjIzIPRGx
mjXPeKfWh9BrFb2Ql5C5JrSdIGZ8PZ/NoKWkmP55Nt1D8Qz4mP2PXP66MJkV1VOtS0Wb8n9/x0N6
697L/2p0F+Lv66d428ce6LSLrDcbML/0WHh64TkQsn5+WXBB6FDrOZBSOHKDQdqv0Fe2mo92WlDz
Xnvv64KlrVWTbCycsOPaYsvBN7ievuLGYY/jymZEgeSDoOXp8a4Xs7qt7X/V05Atwc2sKpO67MJA
XQ0vVexmXiyMgLkmztOka8Q6TYgl6WMNwf2FRGN+kfqPHclWQSv7H004lnq1rUTMFk3YKSMyPYLR
LDSu+3IwPDVzScNXfAHO3cQwlQIl6C6I+uw9ZaC7NZzw7gR4uk6HOvEx8YKsknaA45sB8c7ZoXQx
PoS6CS+gR0IWhLF0KOq1AhaDnwlLEmdbVOv8rWKtuiWUsa5BKK9VkpAz286PtU+4MJ88oB9ZPQ1Q
JFhfjx/UdvZUmeihVIGCzmUfJgx0J5Loa8oy7kWxEqLki/2I4ECUp6dN8N1i1PXEufMYlLUO4TpL
y/Y23Im/OvmvVvIVPMTbfjxIHsv4uMHngeSla1K8iIIlEZrC6dOC9BrTswGR+F2R46KwiTksMKsb
tKj+yhV8zg1cHTwLsiMJ4D3jY3SBvE1JaXbFXy2q1LJlTQs4GhVu7IK35flt4iV137B4SHRp24+u
cVbwAhe9PODoZ8c2/uLeo496pbpUj3ONdryEU+InlV2dI0dda6UUPtq42+c8LzTaSQfoc74aDdQd
2E1s1frpffimJYjIWx++Q/41ZzAiSX2rvIOaaW+8a79qNKfw6GjDrfulcvmk/QFoLRibjI9eeoEV
EgWA8qm1PiiXdPL0k/+MUAEMcKN35BJuTbEr4ihEjHrryqwrlIUyaEsbL6PAjelmOj2z9MXpUhtp
kC8QP1FrOs/QLoIevSeXYImmxnJXvGxuTyNR406oqfaDTyOOgGv2j92/gU8qSSB0Ftyqhif1GGDK
i+ip6qpTmY/bG/JM0HoXQVTa+0pOglfOLqQfeCTP1biQHhgEdOLkmbI6uo68IoGP1SL0rBp4XfPi
bXKurXbRqpxGV9Ce+eXqFh7F3SVHV1OGJ369NQNJ3sUBe78EQUJsVLaSny2aRiOIaLL8OhX1dchQ
yCcMXj8vrxCumPd9ow2XWF9Bu6p+01bhd/6/VSBUSZfi2YI8pXaatcQL5hYAxDKKV+9ELTgfzkkX
F94fGgwOEE+PDysAdhBrpoVdv/SHbUzRPviiCNi6A3yGDetiRkF8/UkV8dqnnCEFV4K4L/2ojAa9
CsC5q3uYiBzNcVe6cvobROq7AR9XbGVfXDR6y5GqWm8eTOSyt9IbYCzOxs++IGjaGRSKH60ws04H
nkvTzNc44NzhRxKMBmzQaN1eCk/IO0RFjbwRBmtHufqe8Uz182pOtLgA3HY3qLtSHyYtRAi9mJko
LSVFdCAZ2bYX7MhxjCYkVQvDRU+rM+k50AvAWvLoS+dTqHH7KjJqUAz7/JvBmzR2Ng3/9fjeE2Pe
WkPCyI4ehzhxbk4Qkw40KwgCFVwT87jrvCXGqKLZDYcAh/nhF8X2E0xkRDy5BeUHeo0E+X09tP4L
mxC/opUb4Ydmh0xXLz4GcLXZxn/Ue1LIBhZgEG5LjX1+5o7H8mvGg4aK8FG9ctiSvXeVBtu8BXZM
rwAvb8f7PxXEYtI6uHCuBvs6NK/ns6h1enVtfYg2ZeVnnqbo6DOry3IyWSHEId9pClg+1Niu5K0J
vzYzPMExUkJW7/Qp98B06Ny+g2oarLIwVujhsP4PKtuyD9xTqoY69aT5supTkW6OycpRLDUBZafH
EtX2yXk3+DYnICjHuAa1NDhYJmWe5ZDFNY2JpD/6QZQzE+2DfyzRqZvEWynnR91DhBTS5AU18p5q
Nm/3Ud4VQsxEj01+ELsYV17QfnCw2KbbKNyuk7zrLKq2/kbXnB3lHOa//UYTev0HKw8AWa8oSz9r
d+0QHYFFp7CiHzEfsTDKF2p8p5mYW1EiF8yP30feB+f1DZocoBivyYdXjeay0zLpMk/9Hw5fHNvq
mya166ZMLfRN3eOI7Tlbx6xpDMp2YUgVoRtVJwlgknt9P0Ouw12U8NhqxOvtXJ3UK7X42ypa/2EX
ESa1g1xgB4Sl5L2EdtqBCkIDoMqmjw+S/BCnsU0AH0diUruFXicJuBOmx8yZRfPmT3wi3pemXabR
HNG1+yHfvn1OlM9fP64EhHn5ltY6d6nbeom65qi5aV2rJO6SeGQqMDs4aT50VgDEjL+OkJisRJAQ
seNga5mUD/3atMHAIs+4pOK50yt8iV8WKGnzvmJVcucgprVFhvt2zQbWaHxGlz7xieCNZqHbPg97
hASy6qLT7LwrJAkd6mt683FK/+zONBQVV5IdVQO66YXqoGUOwTzWEiGv0KM/cKL9zX4KCQt1DN3F
uhqgSYoC8dVl1OzgrSCQLgc6nEK3hPifK17/AxOYtY3Z8LtdXH1yyXYYcXj4DfWRmJCcpFr8WRY8
cUFFndinxJoSNFGCLjWv/ZA2SFRI4mNcRT5qeCJkTUMci2/Oy82a5DTHMcz+4d3s8yWTpFNd2Q9w
m1WyV+75DJLBfI1nkoDouasZe/tyZjVlh8zpZKIlDvDNyHpFzo9GE6pznBbMjXLrEafbdIILdRXB
me7J+gQFy+3cKqumkBlTGM6J6FDbzf1E34d72dO62kLVQpp1xZuHFR/IH2wwLT5Q5g61a6O9kgVB
PGvwvR3ccq6KPkPT7xumIfCJog3YI1gRxRTUMd+igETL5HZ3qVtLHWjNcvfaeuWsQDD7D6R5j4H5
Y2ULxx6RJWH2jHNz34RlLNT894Q/8Qe4Lz2yUuY2diHDbbMNm83futezZTJJZCqGarwXm0TNKOgD
ukA7nuBYbeniWgL8UU9ZQ4DQVFIg1aEuIX1eUcZmglUdLOciwpvlXIMnfFi1dlSBEn1FDm0aILfM
mFO1co/QbUN7nM4a9gJw8jf8V7IkkZ4EEndpkCTQiRHLbZJdeYkcpQCqrb2ji/yQ35JInkrzEFPM
dNpNC2kq8Ys3E0Y5/7UJy77/qWmNlZN7PlxL0qmAtAvqDyd2p0QZ4oRH8PC6g5Dqss8ce6gtl9Id
UCScUg8nahKBd5xdnwqWhcsECTX3FvFujcu6Zia4fC0GnVkrjh6xN/XGMk75bAd9KKHSjD1HskAD
Dj9QIFgI9xaSSIih5ODEnjVXAtlRYZExaAvf8GUtxvrz8pwuKLLTKFzmEIWs66uiV1sHjU7SQ9uw
NvmsKEO27AH+EKZWR+hsWTce2ObYBz9WB4OqgizrYSKHy5CLrYf7jIaezodO7ZEvP90Nz98Np7k2
qLgt9nQ9FFNa4P7+/t6gSgnQYBFe04UFtmIugHlg8RWR405AntDQAlyWRKNhSPNdBMwsILdS4evM
Zp9C8aC+PDEYXg7DcuR8Dd0z6ZLgyCP/e1Ur9aR+qR2DioZMR8izQaeqd8uUpKe15VgT6f3yxhme
v0V7ETjAFQxutVBz9+rQJbOtE9C+7HvUuGn7B9iMPrHiwihOdSKrghvFhHXxwfL0pYkdLJ+s5RBH
4L2PaQPVw4BGbH71CTK/qL+GPv/X9u65cS79RDEWN83F5AKRMNdp2lGBy631r22YsI+NNk/NPu1w
zDZHnVBU3ZbeSCxGbKdk9dtBSUuldFviM+gy2yvKRuE5eztC5egQB3NCApEXtHyp5rSpqA3DehAr
oWBgcF9wh86rDt0BATntDA1E62MXMvvErp8axJOEFF3NLGVGF77soPZMxaQf3kSbXKir5CjsgVik
Dt+zRL7fr2xoL50se8xpgY36a5xMNDjztRj7lkey+S7lMK96JTzJwQ3phYzCaxLYikACHz/Uce2W
VIsjo8953js7agPl/Ie+e0hOJtsRzY6bEYa+YTCdcQSOIno/Ii42TRZJaSpHvdgn6TqH+O0xs5rx
rPHOHIER7G+nKq+8QiFkScbcAlQGYZJ7KlNF4KDXvdgsJPnYM6GUifUYsBr8qZLoTSy0V06gVUxc
NliqRAMcnnTWccG9KS5PrCpENdYosS8WSmFlAIJrzPj7PDc0/g+L94K3YZcQzsxh+ThnHmB5xqP4
Wk7nybDV6kSvGJQ8CyIwsBBlkGJRxrc8ssnUH50Q7iXmoQRCxfzn4QVPiaKjbXXXH0nIzymXTq4D
Wg2n+SooAMbVVq+9AVYktpfEZo9970jFPhccgRA8a7Spog/nhhvWjdBA6BQV51IeafGA1+X//iY1
e5kn9UHyN/hkvUmCJ7RnKIZSngXg5WNONBxTyRGJEugDLPdlCi9uoOOcIICDCAmZc9MpLoj+ml5D
f177C1nH32hCkvNdpxcwbQFse3RJRz0GDNa3aUdc2YTl0OMAlMdOYOkrzGUZBMD2H+55aUV2Khnp
wpwXEm8MqGFnFVCSAnCcDTNgugjhqONObOvai+4a23+aPlXV/qMw/S4nLcHkjJYumyWHlCrINe8D
tP8es7yJrSY2sFzwQZPJp3nuzTavJsvkNcay/ZyNCjQZMfF1wJy+Km3djxwge/TfbWov5sA5U9QU
yACo4WyRm8wcCaG4hO/1ZqjctsdCkRvUjpbwVrpCWBt6hhIXuoslUDpqXMXRlKLGLn9+Gg7JSTDi
6LlVR7v9tjH4JBfAKfXySxpmzA7/z/6WEIypvnF+wKhNNuMiI02jDTVRwPNOyTdxbzEUMkGiAkDR
wo0JzLYvik+2QkyUGGrb22kKvgoSoZScCFKTQlHqhRET22VFqNjz+MMm/LHgEdGSG+X/qVKMbgHZ
nsyAULFntVLQogLbIulOnfWYwaepxI8iUpqQxOXJXYJ9EZ6CkwETHGGF/A90h3Uk7y+2M626R5pl
wyoj92EqUM7J47u6dWDigXG+SUH5hU6p8d86/JLUHXb9ilJpfleDbQB49tLoKNHMY8SJwBY28iwT
w7n1L80/EgeGuIU/hnDHNjLai0h3xdVR8azR+eQjwPFajk/ncOTyXJpoYFIn7xl+d+g9T3XmFZlM
rvxjfxdcc4FFs5L4Euq0RuMSLKY9VnoUZqrmIi8Xb41+fMPcC6GBdBS25uRk7FflcF7/U2dbIXE6
Ihb33EvnQsuXYBza6c9a/O5x19W/KeR4UIuf6qlBpacQA7XN5ODr7tvS8O/xASb6jVBTj9K9qYLq
CX8NzVXPq4+9Zk1Fg/fRBaR7LfB7MmG+D2Qb/J1365hWMXgXaO/sLa0ym0w4bLXMI7wvqupOThjQ
e7iJeLXFs5n3IAuSxEzvKVrETAdM1C5N5gt+YQgj3h3OcVmm1IpDFgo/W6NS7L7HRvkJ28kfg3ju
DKz0q3VSTVu7IXrAsHAhU8iZPQpljy2rkjY6lS4kD4CICt1wWf12Kw3mhrdQwLWHC/PpAjOzAwSV
RxyOwE2iFzpUqnnb3KPOKXDTNCxank/mPeZbMNELQE6E6FQvMxSuaikLslLXMITKR0la7c2aaBys
bbfyxkbyaZDBzkjit5fUDEt2K7rfOVj7910ThodYIJlZnIa0vSKvB7yumVJ8vbFwYc60xC0BXZX9
PRxekkyuPqmT7oZoGUztFq0KkAlpsiH4SooTb5E25w4bWYVWL+BrEiN9jo/W8yQ4aI42kTCTJWAz
vfN9dMFHGeL+T6BvkMGZSef2cRlg7U/tGX+LSMTrC+J5xUx0WzF5SnqOoMbpbViN9oldn0+UCjAM
lJ+SFvAgF9/TaHrA7sj3w/uX5NJlBASY1M77NISlK6j7EYxCuESEDugRk2APZwiTM6dotsA0rRDL
nQP3Z1+l9LfUXMiGG7Lhpl0nvxv8u75pmbQv9yDusBSFCvFKK64jmUTOWyo/fX0hVgDfHDgDJdBX
jpmiX95+MS1ecj/QDYL8EZAls7oEmCg+SykP7dCn9ReaLgX/GVaCKbrcLbixmuqLs7KZktxF3qtt
hs6jBE+ZUIYcdjCry0qCpJ2urmOK2qsprhEQnLeCuwP/dSL1ZnYOUxrGbItF1d4iTHRyBCrspLXR
nFE3klw1T6ktLUQRbLA1KYVGxQtSYf4njyN9OHb6uh38P+5fHzL+OmYct0/k8hYHBSdKKZU525iw
5Zth5tXDARDm3rwD4uyuH+oRZuov7A3c92YWNvNSwacUDp1MmwNA1cfhNAnRmqZmVb8i/dHLjSS4
CxmRVJCAQA51oJvr4XzqRiZvA8VV+VrcdOQbzbilu0Yzsdk+1PBo6VkLX5gzSsd1+ZRnTj63LNBZ
WyQ84CNmJyn/gTLLM39AdD4WEgEjzE/YzhHvnrN1puRYetuXyN9c4ZBK87oldGrP2SSYyW0IzEHN
Ip0ObG/Oor23bv+TMl1cQE7HyZZeLPoFGv6nu8AvQDfVY1BYFBD57C+ViBVu2ZlTUzFZNyb6oazS
dVogc5YgsQSoEAWWE/o5ZBB2DB5FRNvva52jqd/EY67dDIYAzBwebnHWaG/WcTt0aMNSduaRq21E
uGKCmDEu3qkfhJh1EW9ZFXVx3xA4QlCXWE/IglTmUuSt+Lz67Ck8akVOIO++0Kguh94MTgXi2tOl
Ac5XdtKa5R1sMcs77ilf0a1eryHdnxIOcm0Qh1GSyxmzmNbRER8UjGYzaPoX69wfg5YOjS8DnP3r
PZ3xW4dSLZR+xLbF4BQv43AG8qzWXFfhWcWvZXnCOfRe8spenRDqy+/J58zDaZ1TKYV6oG5o57l+
KORtXJIT5bvOgQj472Sakixmlem0bBp86iQKF0KgH0q7JT/2iQ91bd1Yd+Wn/gjLq9lGx1ovp/XX
AcFChkXogJeg3+iQZAK9yhJesvflUbsfU+Dyk5TY61DJtcgN8eqNliomX9Yzv+0W9tSaEYf16Y73
V2z0btMjuEe4FAuc4vyRpGp3DCPw/pehZTDW1PUBDZ4GTW104fp3opj2uSazevlL+dkTd2RpjlJs
4QxrjcMkt4X8f5zjVhJO6m1x7Hh6AHfDv78PrRuR/iUhSuNjn8VoRnPinfQSAPHO7iiCUkbU6Vlm
ThGsIU9WfVMnVGyv5ejYYsY6ut4Y9kpCGv22CV4S3uzn8wV8YJGX0xm83WBHrwJ5gDwQNWgCPI6p
KiOH4nTKo0tNAGafd9aPGFxxfwBVwdMtgqO25Qsco49xXUm5YP9mFj0bIc5p9ZQ7brNE23EsGbhI
6SiFT1gX91ZqYjzyLUAk3n83XjEBImNMCxlJa2bwrOljdXc3vc55S5M8nLWrT2hjtCafMjz/mLdE
PUB0yLbldHGSv3IkuBSq7qFC6/x5WguiDQIN1mMufU/uyHpN6D9uKWTdPtWHjx6HCiebKi1tYyoT
EX0bHvf6c6httTnsbAp8d2rQqm17fm+zGojawHCX7rlw7nJ8iCWHOIrvQAZokTyFAmfH5Ko8uDlK
pa6QNxSS+efIPwVxY0fC3JHYagTsyZxfayZVGtN65mZ4V8bjNqQliOvmt5rM1lQ4TJCn9WbIOKoH
MXFIZqy7RvDneVGkdVNDTsxvC7E8LMlBIx1+SWdh69rHdiI8q7+xofOCoEJshko0W0xvLb9+HnA8
bWrla8XEMUz8ghHU6pyno6NSDRgPArXc2NhrHaYS8/xDGmxh+XHioQ6dClNjjRXnqfrW8gI2aSqO
yZ4DOjaunJ1YFtCr6GsFwK/t6wjadX0dq9VXc55ZKPiUEKuWgWOMPZ5dCOwE10Uncpl4K8WJueHq
I6rtWGZ9AgEcePYKeOBi3bLo0xJUnSUpkS3WLUf9gmr/TlyJagng/SQ5Xlp9S1NBEN4SabEhdrrf
UisTsYVYUuj0xBvKwLbkGKIBeJgfwPzrVXIWRhdhYP6Zs+LHHN8beOhzAwP1NYSFmpTyj8s1ka3H
A/CiRIIUQUMn5HFPmXePTuf08A16ho0qcrzC3L6u0w8Zn9G1Zav/DJ7pqntek+FsB3pk3zDGGFLm
B3Ov42EhNfo3ppzzDT26ow2Ikyd83xdBUhVpMjgusW66UjWFETneUI3HbzCx+ICTSx9ocr15bp6t
aiZoFsobdp9HkamuFEEGih40CHaHdhg0nL4Fy9wwN1OZNRU4mltO5ULm9RPys+D72ad87XaU0Ww5
2sGVfo/QnN2avc2MHo5qjslMp+zoqAgd1OtSq3AmYQpKGv169VKKcSAvb+DItep/m7GKcKTMnuWC
Lt8DmfmijEvDYCfgcjCzY93iZ6RS+2NDksAMladVdRSFE8wPn4/1cd1eFi/EbFRwD7b00HlX7O09
res6q9nvJqZ3p5ZAMgPieLI59Sh8z6nuVGZD+sU+08+7U2B7pzVveO1cnG6nrB9PCRDoc5ApvtxF
IO/pOzQ1GHe7DWGcDXqFD48PMVlMfarO7aA0oFcyVOsP6Wh3aTJr5Wz+0tCM1lDKIc2WCc+MXY1c
DjdzUk97Fnz6eZzk2N4jd1DZH2ix6mj9lANd5LfBxfAJt9wxJjCzw34GyBDFbJsdycv5Vpt9tLAi
dsKUWHJSaPoUD6d62m6SnsFBDnavZ0ZqNo3saDD1aD6fELAiuoDc0fArrsv3mU9K4GWjDiFllg+y
Ks4Zc64XA/kSa8a8Kg+ZkuOOK+n6oYLUsmuXb4hs82XRj6JaOHtX/sk1J4XIf56hG2KIFKh8ruo6
JYCLA41HdeKvXxQrfAG7p5KPJWAOLo/Q+a2qh8Y+zpmDUtzUcF5+gB8vw8IKMLGE81hcM2c1Gwu/
IU/dzt6agITzJ8am25TaWx+A2sLSZIF8ZXIJG+mjeHiABTJVQvu8x+0fZzhtRcCJ8OpZddZwikhS
c54ekCwZXkB8Dzqq+DhXCvZO7S3VB5u2OKbKUAQ32TJXQDTrIeHEAmRVq+A1YTRwSZSEJdmbs2DN
bLdzly5h7dxnf9PQEIUrRNYKrq4nEzX4jyKjK+oTeIxON5XQLlfTWCd2PLdWa3qLVlUZfEEfp3Q9
fOZJ+FwJbNm3YIy69FVSuefnAzO/dyuZsS5x2qqi1AmKdfmmBLnjzx7BM3D23F2VxlkIJz2OeMxZ
t54ir+NaDd7nu2srE6vuNHX4/Qa7bYpvKsUpSgsXLe9uh7ua4tmbHozjMu2p1BWscN+jMNg9Hd3B
A52GUcg3M7/iwN0DthuKXpsIWL9ecKLA91BSwsQ4cOBkeRk+Zk/kok/EHoZdzqXkVahr2WAl0QgT
0d8evNY5SX6zUIIpWmMjzCXlQx0ViZybPsxy+QCxz9SnVYkKUqjt4NSn0Fmo3FUCAIzKxxeNN+Ec
X1lMLQroJVGxLwUusqPf5Z0jhzwB2gWD8lUtwo/H2gann6GUDTWX+DqWtvwVpyznm6VaGuX49W3W
/dS+y5/NtgoP4seknYbEOLq/QDcXtwsxRELIyYMLMP9LPW0F5q4I1kosluh56Jm2aylGstWwsv1v
b50RjSKhjUJmt28VtPpBDmlAhn0v2bu2PoCO2tZSfhgKT4G7ZcGU7olJbBQNNqBLx+aaIIASGivL
ZeC1pOGX9ESmK1oQI0qUodzuuJr76RdZuZF33nzB4u0RpmxO+lbsaoILzyCwEQ1S7Ydaxr6kA3p6
oeCZ9ZymBkt7y5jYfxjoZXuRiWGQ+9KI7JbvToTY3Itubd70+JD7R/ogtFgSrKU9N3pqNNAEzQPw
7A/wCKvxQb1EJ5YYQc5dsx242vkydGi1i/H6HHpwq9xoDLrdcAEtOHur7vkTsf97GKbg5LTj2Ul/
M4CQMkuUiZ4j4EzVyCMv2upWeY4xBNu8rvfe+ZolhbxJv+k32hzD1SJXCXaSOf+jaeG8cjj/BvAF
ABqt+XJBklU8OzWAF/4iCtH5S7+MELbpReV7P7rirx/hZtuF1b2hTm5B/ILm/q5g2ES7HS0gpZsO
THoOq5BhNN5l+jzyIWOcJDfeAH1hhXg6FGjl/07oKHxNgNFnuKvNW3/+89Y85rA2gYa4ncecr5qU
9dCJkA0DsJ8zPKHMnpt6swVSMCXNMSx/O/KxqAr3JzjsSU3cQNfW+sazegaZTGHoON4Qj/gQR2z6
ps8lcMI2RmFk9wLwkAlfpl7C3gdKisF5iq162eUReZumIL+YQPg8CM+6CCM6jkUzp+SMaMIp2sYV
fcXOmmYxGHzRkR+mSs+RkZOj0UI6+5fnDKK8/gdLn4PyyiZM8r/UIeve2Mt0VI10TARlQc6AAz8k
K+MqW1a0v3+NuWG8i1ZrlGAlXM6wehFOr7DlBomxrdBcVKO76rcL0+L/DiwTR8HYlEahvDZRTx6b
eiKnZqJczVp7X6oKEW/qG1DM/lQjF+fxpjp8Q8g/iR2cVzcmg/qS7wGY0+BlXdrOclGRq0UaYnuU
vcUnaCUKMKIG/QtHBnbgfoSXTnG1AgyGB2YheniEC8NrGA+brXvN0aHA0n+bp6wS7zZXVv82qUql
02Ng4iCnAqieJbQ/t8Cp8uFnICZf23gfnilJpXLQjKJtZrdaBFskBAHFmxJo2WcV9T6D3hOt7KKU
Ec8QLyxJ/sbBJF+FRihbn5YSxWS5RetAOjvRKeVYYpKOvLI8sBGLsUdxjC7dmuovnD+tjxv5JDv1
DxKsS3TKHncPZuSUQmvaKDO5IP6cQXS5mw/SkYG6UZV0Qd0n+4/W7lhXGzN4CdkgDoFe+pYvlqQe
EyjXkzBvc0Pn0FQFAyB9Vl/YBdd0sXiWsJZxFxCFIRm10Mc+8XwEhENqHvC66laSNQv5ehkiDF9N
9R6hR7WC82lQvOFu+aceiXelltD+31iWa+hnUkI9w6092Bv1/8LHpiW0Mt9otNcUg2SlbDeZS/iQ
UUeoYQ0wEKzomhQG6BmJYWYcBKc7NYWCXvn9mTxH8vkYS4M0sIJB2Cv5Ilz2cRMzPaeq36ACm9OD
mN7StW5z+s0LjeVmdh0u5QBq47QLaMmeqdgAgpGlC8T6zVhgWImHWTLdDUAevlgYNvV65B0Wpbui
F5zzW+ZiGh9MeMJ7uJX0MZ93t5e7KRMrUglOvlQQSSn4CYJ+fL3jruGZ/6kIHfHabL3BoQMyNPt6
Rx8x2bWz6aFfDXCyFqpfE0g0eVwriM4xntVWH2/Jui/D8qpKx5SPZNA2jju3+6fPqHg5looSbhG3
DkiVS4Gyh1W3GSfzQoQI1lPXeAIZF4UpsPDwqoWRcRABAXE6W0m5/I2nXWifseZuWXlIoIMxWQSC
vU09q2iDDOQc2JUFN0pN1msG++mHJShQEFUVGyByupuqlv4FYwS2im7bi/simZkr6URpXospavia
u6uu1vPXM6wwc8qNd9r1SQMDN1xotbKuDdjCYXsYyc+eZ07+eE8nC3jhJzQWA3wD3uWGW8OPsg9b
2K7c6AZo0VPlGyOsaji7nPffElv94LEllHayV1jkxyERZN+fsX6TSlKdGEw+xMGHmXUEV2U6Wh7h
txxeubWktJF+Ek4RUAEVJEnTmJcLnOJ2mB5RaN9wRDEx+0CRMtEW5xLFAIMmdc6+QxnIzwXBP3IF
gmex21n5ITImrnTtYMPMSewGt2O2aJvLvvZchzQpG56EVnw+Dxyr7PHy4wRHWpdI7Y9PHV24BYb9
MEp+x8Tjx3j/MyyhTsQfJ48Xo58R2Vq1ndgqLZCEd60NjiS3mlC2FM75NK13QoJIEHbi4ID+9n2x
tVqYrdexINOmlEJIzvV+pNFjAgzXxG1j5gDWXoqXy6n9b2TAVYXX2SyWBbTpzugMQlf2M2gs9XzQ
wn/YcYnn9nuaWiNzLz0F3iIgmXak4yZtnqO7CF3Ig6vY86bcstDZdyEUyB3RQ3Y5BBhVGUrarNJD
NzY/7clQrqhXSOXYoE15xa+i988Q4CIagWObvYJw0/tHVOr3phcVY0dixXcwyKyjKKMEwYLLWPV/
tu6U/KdFpCMpeXZzw9WM7Ym/0T5X+KGpV6H6GA1HeLz0+DyTSib2WR1iPuFcbFWHChJGpJU6G7lY
rtPPKEPWJjbRdJbKzJ5FtHUlQ4roUBt6JB6Y8G3RkVx84uFgrE9Va/Lm7F43i2ZuV/wUqWT0zObz
wWLHm2UrLqTPoNfiSgVnpnqj6Ly2Gr5v+GettU6jvRcOyKS6yGGwz69tnFaNjktElz5lm09mwA1h
ncnjKKJX6VebBZwOdiJ8HVPE5rPFtYK9aiygkrQn+Cr2I1juELYNgdb28LYcLltMyhNs4s6CeUHk
isfU/vIlq8a2VL+SqQUiDUyRscW6rTPFVaT0C3TJ+1LPSYgR02V3uBg97rCVm9vm9KtPtSr7pbCG
XtokyaNPxdmRm3QvKuZC71V4E3FGfA1zxGWP3+fokRoV1PHuJiyiC/JiSpEGrVvdDDOhdUs179GA
x+yNWm3qWVJQq73zU2t2dUkczBWBAh79sHV9kbeVBqW94W9hzUuv6tflV/Y8EnMbteTmqkuSXQcJ
x+gi2UOWwdDL9zm/Bz8muE/3JHB3V8+xC5MCMPb0KThc8kev8+g3xgO1LA1lEE84SMykj7ml52Dx
cGNbDPzbUV6M0/vTGuccAg0sPqO7T799BVULNuioDRwixGGAyKRPZ0rvGdZd4Z2SScojUVEu3hLO
2TEOrDDDHwkOhts+9OQDdG505t+PML5rDwRRRCS2kBM4H8qaoh1oEv9gUtyLNCw3/6+bJ9Q1zfiv
ASCoYlmifbXWcZKOhCrN0KOdbXqThskebktmiWq/7DSzSz4CATFX8GdrF+tgorxAreHAplpgBSAp
4TUE8JcitfGUQA6NJ8KgGbbAbXT4AuNY1Opuv360HxMd1pcUB2t/MPagkL9OZdtBvFjnMWBrKq4N
k5qo2KKu2r4tKdmnknmj/yaRffKKB0KvDbJc1j0O8oSRj+5BsOrFZfKSkVWVu4wQlrwL/v4ocIzT
+QwAvWSpnPvCFJT4ufX+1YDgQm8jQ02BHrnh7i0uTBYh8gGIWdLVk2qJJVFSDs6bNgE7XpY8THm6
AlhhC6KiIlPLKaUTuIk+fiSQ6kaBNPjhfNoDGLEk8+xSX/Bk7sqLuy6oOUW5WAfEz049WcMJh7WD
koknKpVp/x+LkKQTakDNQkgLZNxcop5WkoPRl2JlQnLgvjhxP8cNXvpnXj00viGzWUiqkZf17xZh
HuyW2gEEMR9hH5OqkmLVANP2MnJxHfrsU4r6huh70oTS5U47TlIYWwTJcPIIuhvmC/tQAHtMzWzH
hvJpAuB2kQLpfakKPU5qDD8O5rdMFHymQU3z7gHBx0mW2VS3dRfatZkIkqnkFprzu01JWNYvTy+U
O6G4pyz8j5U03TZSXlyEYE/e0Kcd7dlJL9/9YM5/aLI0Q6b5oiIMmvuQ9nwibApYNziTfJUBgJZY
08FoaIT72vq0lRZjmtgkqqNZRhD7jk/bb3sTwtycgnDHKL1VPpUpcrS6kCIjOgOHcuscxARlnsmH
rt4/+OSkXSOvubeU/Fj/ow5q4Nif94nXk+qXwu9szpKDj0m11N1kPEc7D/lL90IIvi+TOVB6Yx8S
8bCuWwQAfGcoD58KNsh85Vq0JD+QJH3qiTHOAHmjO8Ze71x+VEn6Lvrmppc+PKDQWZsXS+k1RnZE
goD9+zDaeTNOF4y96geIJw5UN4+IYEjAAYCfZl7GAZ8c+RPfiPIWQZThsgr2VXH0t/o/oE8m7FfB
Wg1wc8kIXRaaEKJxZyGqV2VOsQVI4W3unYQuYpSFTl0YuBIXFEVSwstU1NCHAjG4y9fcLY+nLc5c
k3QgnIczF/7RAdI2pcpbRHS5X+gxqF0umbYZ3sU+lmU+7BuxEC1nx4NEOklK/J6etRgyHn4DaSrT
O/z+Zg9GPR7AFoWVj5LNVjPwuoBv+rQu8bScE/CJKXkhU3UUuJvNjZ0VFpyXWVjR1SJzmsj/1L7q
EUpBLcTSB6vf53UtaH+ari5l5yhYmwcv1zfaVd2UsZu1weNcx97hahFxAFUEy8KN0/czu+QPVHwx
0Y2b1FH2d/0Lqw4RIwNYdRND5b2R/rfZK83pDLsksgGVLk9lZ3q79J5Xgdkg0CH0hCRthywFzsym
0/6SHaeYIxVbnyrS2E5nszJVAhzG5sEYyvLwUEMAK5XdTH52HUVDFKrUhHqefjWniJueGrcfczs4
HS8Y85a1Mc6Xzw4IQ/Jhg/pQ4T4elO+HwfbacK6YKEU4XNZCz5zlIT6heMTs3qIKci5Csnp00QeH
Y6MZWhkH0bY5ME65PUSKQH5hBEPBGSzHB4YTYoIsKNFk7HoVfXDbYP28RrjZeLNKfojKo0NUhaus
er0YMts/Tlkd74rlYkMabGQ3+KZtWzvwCJZodrVw5ZgdJpVc/+pnD3ed5ZETEoi5Bory3XceG068
n6M1Dv+MDHvprWsz2Lj8Da51YQcsEBGTivMa5lw3gqFHjZmfcjtay/+6ZjLtxymih9zSovXtb02G
PQ9Scb8Vs8otcCsWS6q0EDWH8UwVPtkIr0y+85jLKuQU1WhnMNrYJfTAgTjbkV+fD2U8kQ71eyqg
YURLBFz79LxYLVbEQ9ZhhVNF/RG5jDfOcmclrZ/4s9O3zA1qt39B6QOYMHNMFSV+gR34UXHwkzIN
XXUsArS6CvnU2Jd+VOw0jdLnRh//o8jSI8quINQM0f94KqwgugfuAvdkFKRZ1Z3VUoNiJHY+nJe2
G0ehQRdHWDZMza5vK5zqbBZT68LIUt0p7Q9mTgjqGWhqqRdyLOWQDP9y6DVcEP3/wlpFI80AEa8e
cQj/8UYJ60/BZIpO85+K3c8Zc/iRYxEI9BoDCNrZ1e85il+UanxSeeDdvYj5qZ7A2fTSE20X7m2v
TnsvmZO57b0SqvGGhDmaFJLYpuZFLzYUIPaq8/M8+oRmEAGaYU9gGlTyHh21edWHQsXN3MpVIhxd
owp9gLm3D4SWjK2/RW/ctPANDhnFdFrxS24YfwOE5k6LmwK9ED0c1M/H1T9clREQIZfiNNh5DBrG
aWE1ORA8HxL544rI0bl7ePJnIyCebhKVe8mp/hcqzctDCNsNjNmhqnCv5bdopJZuPj8MtV0vHl89
MSlFGMCgvgNV9PkY8imHwq4cghN5vgcaeZ2LzlLtxMSyxTvUIdRYftRhPfTVTI0ahT7kHXIOzYRn
q1X8LOEhfA8XqDwvCcUCmnOfl5HY5eBK/EiEALYEs3HgOor2U5TxMMPG0j9JV8HNJktwQvkX0UeX
8OOKiCmbUZE9dQMgbmsvkybMH1CReHNx9fFHiEkBTSdv1WDnGnlazCvWDGZllOheVAbZ9z6Gj1G8
5biLTluxE2Y1bTJahJ+2GBGcTnFV33codYrkpf+Jyd1GpURRVZ3tnlieCjZt20PZTgay0D3vddBN
l8UG7ncseHE5fcNIjrqWv4eUbz/o30evL+IfVyjKfb9KXKCzFYqY5IhiVKwPTBfIGlox9CbqfgKD
s0zximdo0qKFG/5N/WPlcv+gV0wc52t+Kzhv3e8vR3eeDZ6p4yJfM4I2uICeudEnMD+HkQklrE7B
tXgssmhSKRqd8QJKtaDYmoud9A/Wn/cgn2qEawdRd4TwnijzRwV+XfUJgOqWGJNLP5upgjn10QEr
kD7P+IxL17XLcQYBJuetxfKgIfeNhHDlisHWPHbRec+nDXsd2neLPBi6I9B90wX1qWwnW3wOhDSn
Ik4wNGdAW2GpZSegHCq1fV4dTecXcCvQg2R8nB1Fuwl1NbZB1HQGG1dATTfB1/SaYeWzJd/8AzAc
nPlM4nwsp0KgHCab+YCLA8oLw6JnoQEsujtGEDasHdvY5/JgT6ztkR2KO3vGlVSNbRFccfRAP1zD
//Sm/Qw46Dfsxwz4IPN2MH5VHe8QMSgjmGfjzj8h/xYfnSDWEZk+namHdpDL18kpvP7OwbRa3CGt
DELgJE2JWU+dGH46nysMCGB6pHjxdFFJXIYep6DNw3TBXjdXCGssL0IFiGV1YkIb16rbuAxyEi/l
KC2ueJYov17jdmshBz6Ppx12jLaMeA6yUv+SKZsYcuF56sxKvBVci+Z9acNbKVYONO7m2h2a/G6Q
dFyWSnZ9A2N4E7aVPfDevvSur6AzZVe4KXWmnFli49eL1Sy7DTocDw813wBg6NgKwmn8SPLIGQvp
MCTWbbBv3b7jAOmPMkARACMkfDS3hiK6xQ2VcWRlyfd83S7HCnYTepOM2Lx3vbD7pNDXMeHCz2Dm
w7DVKTAOghXYP5eZFbEop83G8v1/f6nXOXuY1ry4plsIypdj8S7DhA5Cxr/yzAqDZBIJBzHhBgyz
cHi8vtytg21SkNtE4OYUh/oMEjr7tHBTHXqzZgI6RmEIbCgUrg9DXG1EI3LeRfAkX+uW3qPuJWIq
HgcJ7q2qjEWbQGrNBYV3zXkcnPPQGaKdUcltx4ksmu/HSnunHO+cRw9nP9GUx3dSh44+gUEybxni
OhkrZWUfm9I6lz5XZ8v32XY0mrqYyycez22h+jjzSvEfyGyVDYPJc0Iv2pRrDodClQNeZo5bU6s0
MHahBe2gOeVg6M1XGZiucTsyhBZXeRtjA06g0tKIH7txoeIcvNs/Nwl3rENR94CnJxTZSrT2tucW
fhe69mMDhv8ZdUFBKNtCTMsKEz96dI54UrG4URzQ0l6eQqPzQWTepPk4XPHq3zC1PwurstU7nu/1
dfaCbNDgu/YWP+twQktPuhZwAj29ePhvyOSVuHVye2IYr/VKlmq9zoAen0hR/KQ0KyrGfOGGZNLe
jUe1+/jCLaE8mUyZfWRhE4KpBFX1UCFwNaWEkkaDKCwCENkTq3bwg5QS6slA/pv5AX4+H6TmZ4HU
qN4R3Bc6J14+2j2rWBEOeCODywBZhUk58w2X7iPHj4jJ82B8KkGB2WG89eeLUJx6U/xEFdqxycbA
3mYsTQZoT471L1BgSUQBW8v+nrqI1l7UivZs6CrmsEv9qu0OIrcDfJkKVV4UEmta2rcyPyJ/9SZa
yrswxApRk+d+gTsaMo6PvT38XaDFUHDf/dTRzChqL5M7ikhv22jj+48fML9+in4NlXcW1q+Ek++f
hqQXKYAWxGYKSRjzlKKRqdsPPEZ7f9T95qRTYTcUC7wvW2DPlLL5y3WrEkh5sNK/twjTG9thI7vj
SwzGbIXaZfjzZMOFwZ1AaUgFfisIAgH5kIsgAtH18PXsC9v2wjD/xa2g8FH+w3SlSuz7uuW6RGGf
MiKhEeDVUmhQ4fIeyUE2q6O3NX+XjvlJq9AqCm9+Yok6Q35iJhuFrFIeWxsZu4ZvBaU283xKctj3
AT4qfiUKpYKpcf5b/hlkrZQnUNBT5bnp63IjRiykZOQB+WCSIr6QE6pdrvIQZTByAyTjmh9gFlO+
jfVbuu4PBFTrOCq6UM1X/rLTOuOtrrBILrPCSDVnIzcYjUrY5CDjyxgpjsZKOxNvMAAXLfMViVqB
OuEVdLCfvrrtdkg1I2F019OlYRzhqS/aw5tXBbXxz9d/vjuGpoFkDOZHQKybviyoDsdvfW9uNTSX
yIJq0qIGZUfV3HtRbwNOWL3MlK4V14TCt9oegaX661yIyAKJr2iS0CfQ/5m4KlI/RiaagBTTn/BY
V+Gl3+pCmT8WCYkJi8veOzFgOK7wAytk4jv46LsptokncFrAEqGEqDcRJQ6unLHRmR5DjINxIuU4
r23UQtCWqRzeDi+gxLfJ2ylVwqazq5cOgt1y6rpz+5F/SSxfG6UWO64vtaZ7Yc6t/68fjI6kJeIZ
nIX/KXS+hVGsylKdrkAD6N+qUxBLA0GrzzcW6LwDA/G7c5T1zYzVnPEVVw4yU/h34DmfpSfYZREv
gk3eEMluH7syNkujabE3DWzBpdvgKjgjmF4tnK17cOBfb9iTYlyGvOFKPLTROxtnyzHapFfKuoOF
BqfhpJ9jPNGA9kFc6uQ9uLf84UILAkG4uG9kW1//+nMjTWUw2EUqSthjwZiAKSCRWLg1pSERaytl
xTPCwyNs9Jpmk8quIOrW8yI7d6gI1mTMPXj/K2ry85/wrN6gNSzNo6+7Qpe2b3VJH3ry/O1XEb79
S/cdtVg5btrroRKx/oKzJv3GTBWLjJOM8Z6Ve4kOUFJl9f2DWsTDbUPz3kJdFG0EN0V1p/lMD5YI
V9bWNYJlxrnJTk3mZbR6BmeiAos7ZjU5+6xxzW9bQTH/77va2h3hdmNwxqdyFzKgpIwTJ3v7mNB2
G1FC2qHxQpN68gfV5kPhLLk9QsDq8GDQpHB/8ZtClcpn0XKLo3pUVqIfMglzOAWYNynQqA/cTk5Z
ir1+axM4PgE6ZTeLwDPrZ6NDhi5H6jGuqrMvxB+FwLLO4lEtHtz03NfuWgpr7tMsVI9HIVvlQ3Zi
inZtDn+lTWwUcb0K44KEtuL+JNz2VHNlK7sWj2jC9vfm5nP3He2N+9rsfZr3imfSDG9zq/YoN0wO
CyttTPL32eWma4RDXfi9j4lZ2Wwik2gRNtivOWhD7n9NwIqc3gCZgoptQnYDLUtHPh58auEU97rM
kdJ8FRnbzE0gjnKqBAFRN0FgKuM9+YybhQYBfdiOk/H+gT6HYaO+MCgRWl2KDDIA49amFK2teHex
eJNQ5q0/DxhTxBX8tg3v+j++X5+dqBMtmQdMDJx2oyovLwc1OjFtAIvk01DCOzU4btpizzD0AQHY
dW5EWe5BLPhoubijYxYIO5al3rw6ZDuPaStzd76zoAIwt0/mj46Zy+CVgm650iDQ1yOR12LiwbuC
JDR7ah9r2yEi/v450GVbyeINDNG54au5A7Z27HdMgioyXAiy1rbVUx8Uc0C2EW9L1Aft3pEjurAL
KDhCiq7kUmvg7q4E0Mkr31/pB2gyqg72moPdH1D0tSlkjMcLUa89SoD8pJ8n+yRkUBx18JLGreWm
xkVAILiqJ/b7q22w6vrn1LqCKLw/tAWUHF7lfRhDmcdZ4V9vGA0UpvAva3sxef7U4P+5Z4tirZFw
/XG1cAGeVagHOM3TvIgcxfuMqKTQqHjmSDmKpD+oub1h0hX5TWAVCkBwMLDrdHWw/RKJ1bG48wxX
MpyLTRlX7sqTLkEdFD6Z34HMJMEl8wg5uy2g+qosGCQ+VVweFMW2VIHgpKRrzpCLq3PcmaOoujAD
IIkYb8pP9a63axuKaWFYYcdGDny6URChgjKOElyieVgAkCkiipnz0d/Ll5YcU+lwa3CDVw45Ow0e
e1j9U/T/MtMzD58gvhKN1PFV+QuUzXnuqlgHJAAEWDR3NytI7AluvcaoYz40GJe9yNTiK8qHvc2O
V4WV66pq69ni6Jkp2lEaREMNKiBxm9+yui1E6QtJITtGbIkvTIo7WvOiq6sRp1orV64N6DOgTW9z
0I4rkbrgItiwWfrtpHySzpRxB28Cv3ZT8cZh31R4f5+4bS3eaKDMSioQ1VnBv8toajjK2OljQXJ4
GU0yGE/bubVlbuctT8wWLBJzK3ZONcVJ6BIguxsQRpKw5mgIT1SLjsAw1yt+sHYnNB+eFvJwkOI3
wtCEpPPhpH78z8P6UIiZfR9Z4ADeAFSnrSJTECntwzjQlV4rAULWqTnXxsc1AZjaKd8mEq4rLxVK
FvRUBmlb3IidO9hiaky5BpuhhAK91Xwegl2ZOULM+qBN83+86hhfWkwOV8nkZP5jj5s6ci4O0Fe1
cAM5F+ZeBremymr/1z0sqonT2oEzhfNiTMWp7Y6+iUYTtGc3mRz1tOp0RC/gzsDT4kh4RQdlATKU
g6gm5dNAqiE3MYrdGAuonFuzdLABucXP/lXzP1/v8MpPFSBiUrocXsmPND6wkZZxtlp9eitdUKAX
oZfZJMy26Q9Np9OLuaTT7PxZyyxikHW4sItybvXPFANgy1wGebgUBeVwX8PsJb0iYKSpecjeUeMu
NUebVq+jY40gBffs5khO8e+OjlAwVeVZu0CPF3/oQ/3g2M7xYg8VgWNTO5uyIYLO9qirwKbMuZfX
qUO/rTTHIUHWxuodCkQU9UQHNJqGCFWxcCmVY7JcdpGkmbAXvOFwOcxPObHzTkB7irfbLfAsyqa/
nHyQ60hnqwO9V+kxS0oqRuPtD4/vroltLvZqt9iJHtyoNKViDdSsO6kkSHMzYxOF5H1ud8rk49p9
0Zeofk7odKe0fWYsYbVtq3A6oFUMib91d998TfTDYHLPT5Uomagu9UhKfA4G+sBIDyuP1zlCqhG9
vzah4NB0ZD9uG8pkeOX+/CQBFibShVHo1aNS0gQ1872SLNWppNb2BN7I3UMu2h74CVCy+rqPJYzy
ruV93HmG0Mi8gaHOmOuxF5Z2ggyGBhonBqLXAj9ymh9qi78uwGd7q79g1qV3jXe2L3Xxf17VytLY
MjecjKbHgvNarw8uYHDTQSySml0B03uGzWGFqBLbpiawV4XiiI7WcBxKfNN14bqlx+F78m3qu3dd
E3moDEnEOAdr1kX4spdvTumaE3BeP4gi/t/s97rds5cscCb1F09Wdu4UhDcU7r2BsUH2cufStbub
4uRMhjigxrhJk+v49AIyE8A0tSRi+YvkoVMrS9i7q5u7evH06Kn73elcs8yP5TrwJhPJcP5KpfYl
wFjrJWVNjJj1uJ81MK59jdqfi1oVZHRhpPkhxWHgTCnkfS2qe6F67/h807tFR5W0mrToS+1DtapC
7LN+Me4PelTsFcUW60SunMrY+xf9dNWau44s9K4lXLvERkLRjSoA357wP2RCslo3noJdEArFXiZC
ss2aR7DH9a1RTBMOFM0cW/FWitjF/LswEDgvNIY6hU4gUeBeBY31ql1rc4ZHSazGJZQ4v9zGxNU2
5hUMADcD1QuDrENBy51RJarw9QvFPEh2xRpvZ0a/kv48t5xtdrDCUOmV0k9hlyAAfciH9DWp0hAw
cquvPtPnzTM6h7/ZTaL8RzMMBxnBoh7joy96YkEGqJkWkHtOERtcRjBz0YYMi1gxhq13xsfABJXL
O94WeLis+DUquUKQDW+Cx55B/ef5l8WL5ilI136G1pMjFBakfE5/YXAkBA8MWONHbzGKqkkf6G51
tJxQ72NzUWEi/+ilreUrL24NO9/IsKHLd/3QyFAJ/JQQS3MMUzmSmHr8o5jGXXdM92zxkYP+EybA
2o9New5kQ8QperSqxA24GJb1vdWia3hOxWceD39YnbMzAEW2x0W9xXIRtQf4BmB4znGkuSFd3s02
gS5AP7fsh3IuQJUzpLQMmwgnW7MvuHb7y7cw21HIMPU/7Em77CbPKYfuJ3glfx6tgJL08vpYj84F
DSMb5894BswtJm6nzH3cylUWvhPdR06z9nlOcpyVYrZfqtlSGMu0W3OwJrn68w2yGzaeMqFXWrPO
6srkhaw0Bj9jYdBEHn9RTXnbdQ5e6GdnmD+DzZlZvlCaqUoH39u8U6cL3dX52Ft+KCEBt23NWEn1
N+PILY0xI5yj+uBLAeePyIxCZkABdknY5wsi71rMxEk1+3qHusZCkof+e53QoJzkG20bzvvK4Hwf
mvaQQioaXcF8OXcLuM/e0sTRyfCicFIHMvmURRqM8jqRcW7jhK+6QICj3IpTBTIzr/YQ9wLR8IXp
pN+cyZZxpdnS096X2mFeLTdRXhOfFLyN1Nvybo6o9dWPVy25cwjufrkMQAhSvZMHCN/QGanc7ItQ
iHTfS+fA5zgtyYGwMBJ/JQ8fmGpOir9yCUpLb8eU/ppOsIO7O8FSrY7Y1Pz9eWGgUlA95GNOVvUH
GGcE3z6KXXyH04aTbmXEOhuonb5JpYRxTxE2G27oiU7+xkVQj8xEnPX0k4msSDlzvJcmIVJ5MFuQ
ZqZKGjNgOh8pkDOe8Y687Sm54OIBjKB+i5cFa01PqJTkn8wn51yhdHHDht5bjUBjxImZJVNq7TIN
GT00yQf1nv7q7qnffQeHMv82tYcTDPPPHWftY2za7Zc2g2aiucsmzU86JycDt9aBmZr8RtVDaLqV
Pzan3GBuVkCkyNTx2zzYOQu+EWF84exxzS/XNbnHbeQula4iqLq4g5J8JJi422hCpJXI07kp+7+h
x072hcBjb1m9Li5I5avYpqL8vhvo/ZLGebxDLSRJqCRp5IhJwLODpmZog7+cEggRCCc83ehpwhv0
MKOE7dlpeSeZc1P3eTYgZjiP80Acvaf1xuqiCwkcGEMQQ8vmhl5G64AkccuuwVhR3HvCVDBwouol
1EhgN20nMqK7s68o03Xc4POdN9IogqZRrgyKdV5cGaGoTiYW9nxLQkCDjT7Bj7QWPgpJ+oop91hz
U2nvMeR2z+J3D4C8xP3MgZe0gclkMzY9bvOdAzDSBQqAiYTqwa3oWqr6KsW3se2aYO1neejxtJhZ
BmFKapiK0iYYJCPMIat1PbvEWTPrk0rVXl0UsQNocImGBpSBxiXpeDI408Zk9gWDjsRoJMy+7yAu
LjuiesrmRlNmC1o8Ptu4rLag2L23mxQfeBba8NLh9XfKfkQhS2GSE3E2YYlawuBc5oH2KvD18Mws
kurQa0BL9NXn2SseT1DnAHv2AyN9Bwb/c/nhrEtS7mKyX65UCbGBZp2lDeiJ0AsmiJRl/Z7pejXU
vLOBMPIYDrvCXL01OyRQN2zvmqVTykBBkwAhZCZgFAw0TkmDPbdNYMm3a87A8vHfjJAHB/4cJLOE
nfSlmmg6X0nrEzNpncLMwoA9R0GKLI6shfofjLor2NcipSkqbR6XDKb073JqyhbXuB5DA1qCrvV8
f/cw3VY4tyy62dkK1v4/JvZ0L0FzVc0XOkzgbZySWAvkIVW0KzRXIt8ZQcwZFbJH4OVJCfkOQnXC
xcMPwfXkyYatdeFQC9BIRzi2U/MxlPVexNLN02K1nROcziw5GEekMlZRQtiwFEm0yowMHoyAOuWO
Wmlp9obHj0UWRpk8K56sggL70GB647QXzT95XcY4B5ctXJSiXGXprf7XmodR2M5c52oQMk7HE+Xi
V+ZZ3gUmZDhgU+AelnNqTHrsEELjAjcG50/KoVkhMEdxMhZGUtTH7SSi3UcQaRB/xRWQ69+qqVPx
E00eE84OMz2ra4pwBBSxd4XGkmjGuiT6dw8WS+bH4/+Ju8Bi2pZzMG/p06myooF8s0HHBu2EdTFw
eruN59foNz+1UZuTFeZDWZr/W2mMuwOKwAe83NAL09q7pIm7lL3UA0PWqfyQLlvW03BlSzlVmMe7
1bxyLP13SDnvXO016K3y4D/lCmSIN9uhyWar3vzQvxQdvPJKv4kLcklLP9Fiq7STJkiURmgy6qCp
JdTIXD1sP3tdhdiArTkygP6DfyyF/9qUDfYJC4GaSVd8r0vAaQcjJ7gCBuhEiTZ3+XA4Hbagrzk8
b2lDkaTyQ2gR25zH6WORAcZP7XlGZsYzoAIhO46FfJXEDMR1ThHDVHcx552xgg134QAmsunoM8lH
ATQH+uWioIVp+vCTLKn+/2tpsBAzROr9C1QL5BK/tJgDtcSbYFesodMLsanIyJB//mwLNaG0dt9O
ooAeX3m3E9WOUerjQUh9ObYhS8ysBK54gLJLfEn4QmuLv22bR5W7yPZ5g66/7rnRJn/AWfA0zmHG
Lx3TJ/oPFNXVylFbfFb4Tz5ikIVUSCaGBqFWhgGaFAYWPudld8qs72pDxIFF7ozx/oUo7Bo6tIgp
Dosd6fYc+HGrdKENRsE3JbuTlcHbfRlBVRlr/VJd8T14//yhB/SZdq+8KRyo9Pfsc52RRVyzIIgu
Jyr5T24bfqWVp4QKiaodOTbwHAB190wbncWhk56sF1S+cvHMwD0G2XQBfh7hKR78uiFtq1Xn0i32
uwEzAETp2wJN3DQLeaQrZnXSahMQyvkJIesX4ID8artzgq2xYWUluPiwiIqMOwARsBdGOs97LE7a
2vqHx/4oMbpgQwr2u4R7QwSA8RbxD2jhjs6/V2oEgTGttc54MMrjWqlLtepDqn129/h9PSyfERI9
8W0j4KufV3EYldKobXGfN6lzl7UWLbQGxgVCev6mSunsRyuH47rqH56CzEPvW/WcCVuqPcDLv3jG
G8DdAorOY1tw7s1gXrg9QNZYconN8IpXzuIOfyFEZ6b4zuF9ddOkzzjoaqKSue03rov4D33Gqu2Q
dw0OTsFQHQtUSglaOM40bMfve3uCEnOTPdoMra+9vjiJ44EvUm/x1PdZ77kJeEICZt/SmlKMCToE
1W5t2hOaHcKos/0f2WDb7bG/qENfo+RB8Brt0R2tMlszzjTkD51T/py5HGLpGaQ+/4RBR7PiOBEp
kojRoegRE6ab52yEdWDtk/0X/ULuSpqm/ycYT+iYevSKx4B78nkSduvB5Ez7aFvIsTc73/v1YNOu
StZAh/6/EKnw3hGu4KEvbLjs8b5OdsyOyKuNNNdfaO+FeCjHojlSYDledPt6UgF28xLRMRyhJrJ9
ROLAHvo2wrjKLVJh1w8vFCaM8TtxX4kopXCuvKShUjjZGQcvK37IUrw2isoqoW3XE7gZv81o7k8i
Oia5kPSbmvCKIMtEy41yEmmGUhcGq7x2AjIBcI0bgGXwuhi+gdTn7BmnLzbtz6CLtnsvmXEkzIJL
aPmCbnY/IA0BiJKA6VYT6hQ3LDLszYSz23HMEjKuAomMAD+1mPVOmPdVdWdy/cCnSqDBH4iQON9f
pympNp2+aIx/W/6X1AnKgG2m5dAcKEECBO7I7B5V4uhmSM6Y/Yhq/wH5m1kMmJE3YiVN5g452Mbc
FgcFIN/aF2xv6MDHzoVvvjWZKN9WycvFL4btRWA946Q3paRrMZGJe6p1Ps/T5qefTI2rWyhUSaMV
Z3HIuskrPEdbAICe6woDgeeIds+VdXwyXc5OmDuTgXJzUJkC7JTbybeet5wCsaH7dovo3ryv+0Wz
9c7OUNpAzpVJ/D2Ko4NwxV9dIPOiXagrXCos4h8BDokAS7I0zj8fOnXiVHq9whK9aoEz7wYivkld
VX4QP8tUemPcSFegOIlvUt+5eygK9qRmwe3j6zJg2VkXvNsclp6JM/v2DTsiNhtofEMJol/6HMz6
nbm2UaQ6J3SHTkZvQ4dmSrW+Ucp7SPvPZadqro1YaOisPinnhDvVpRQDWk0wqplMn0xERuv0dFcO
AKraUu3ZUpIByfsaMEZHBOICXt3nVMaDVbjoanXI1j/YmCjrI55BlDJj1F/kImfOSWqg7PZE9PG2
KZ5ULE9IG9jVAlKjd0St5Id/9IpApGNXXZ2VwyQ7cFF0EAcu8RnN5WXp9bZ3UGOKrCF8oA5/xOX5
UJa61/6lhwP1A//t/xGqpX8ChsZRIGTJ0DJMATmEzl/FMU2pPzL67m2ApE4hGBjPF1xJ9K60h+n6
/kuXLVG/Psuf0DdhTHSfAL/VhTpSfo/m5gPRwMXjZSmXjJoE4mz3YNFK24j2cU0O6jufmnXql703
G7uZMaHcPXudW9KbQ6M45gAK0f9mKzt5FneyIL0rQEq6MkqN3xaUxNOc9Fj+rb98NijmWlZaHOGL
AavpsgGESkCOXV4e4om1OYeOZCzQNA9R4Z1bOEoJqCBdIqjepZQq9gMIFNkyGtcCkjrUx/Y86Nms
fgxTnptZXbB1djC2veUZHfngjCb0Z/oIm+L6ceQHLRitsN6cqF8SBrRvnNwWbSJZRicjDqtPf+Cq
tdUt6U47ZDHWswBtD0IY601FVW7ZDRLVIlJ+PibhY0ZQ6yVMRCURYU9VORetBOftSEw5XNwmvcke
tX2r9Gk+294JuQ3TJdIw7kVE1Z/GvpsRyplQ2Lx8B1Y7XC5oaYPWfrOGyll+aNkmRG//6fHkDu+w
kclaZL879BquF6nq/WpLt8EMzi1rihwQ1Kfa5lZ+uJitYY4nMOv7Z8BuP/nLCv7trUX1DAp+VAsH
CSEfVEwdlgWjHR4RF8bRzBtdhDtK5WyLMXBIpOdu2OUEAszjCSSPmT/NNs7Un+zWM+1Apd+jNQth
rU0StYsEPdgOKzGRE8iaDALCSyAdLhPp3sQF4yGP/MkDUG7uRomcV7hDgDMzb/WMG/u+nsZvAKz5
byWNym4kJ90MTVqGn+Wff9HbPRUNJVVB9mxZIxJuDKSxf816SIRO9nqpDRarqwSzqSfdzkpKIIYq
E/ds0ar1CSnFzC78Bo4KihJBWETIkLMFxujkBEyKHrNUZW7IPhRZwUHYR2EsXtmgADoVhtSyudqZ
rtrAD8yodFSd20RhAtLZtxd5K8/ukCn4JVWrsK2JK8ORxHpWn2H+GlbsCNiyiC66vyvQkPa1bMSo
xUNtvGNPtdOed0eb2ZQfLPuL/yR+RLlYp0s0pp9uA1j8Mg3u/rB4Jr7Map1VYBCIX5cbckFibsyx
nQph0gGDhbd54YvhKvGFLjVj5egHrxnd6LQACPwSkSZgAdtYq33o+rSvzmBNU9b0g6Bapj7UtDze
dbLiBA7qBym7VOqdB0TEi8rOFMKL+07N5ZIpjY2f8m/khGcMeFJMDbB1u4cDjOJfCB5tuTrb96wj
WC5XS6QhHYcvVW5ASuyxL4spBaR/iHy0xazEBUtOxiNyPQDtdxzb2UCWIo6Oz4SNJh6/dd2XJPSi
Ue/CNSToYGx030P+M1bXHCmS59BQa+lJ2XKdjKwtJZKLf3xYE4pjGBeW7eNyp1pm2iIqdbz5gsyp
Lm7IQCr667Y/+n3jwaoixv8uxfBCY+o9ersCRWeQmrDmAYI1OsohQ2KvlliPLuJQ7VZZE9/Ui/74
OBeFlhLRjAG21ofE5BNHwdxxmSBc7CjhOqbjqERA9wPdHMRdpscacq6WfmJB3EL0vgwMVPu1Jexq
3Q35bbsEKQojmLAX3zb5idDt8XbHTm7ocZOM4BMzCbbFeVAIqI4viM36+APRnjRxybYs9dWh37XQ
gYghDebi2FseRmsNFdv5vNwg0mwNChGioXTOR91Qv0HNcd6BvPyLRXV2HuEY+VBVgwnUoxzb6ITD
RxU6njY8McyAM8JyJdA0UPZyHYyJf3yZl0eBp06+mUVQdxkrjarA3NOqSzNDr/ykinTLQPl7er2r
DwvX/23ppCHxESWp3DtwH+cDMSSr9kRlJa3fgmGImKB4GAc7Mt9O500JDSvTaaiyniu/ZfU3eCkJ
6fclJFXkKDoWH5OQNt/nZDB4A8igF2OF1C2Qm/AvRBdmazIxUL+OrDMqWc+tsrKd/528kiXRQ3Ou
FX+0+8y3NLUcO07muWdUJLtQoY8KqBRqhuMi1eZ81PQ98DOF5J2Q2yUyE/EAbVTLgXTmZd+40sbu
CPGLIVnj5aBSrm5FimzuEZsZzwg23phUIICF85/JNRg+sxQ0Ioap14R6P5x/XDp+JnIjn6J9GU6t
V7w1FFsPArrI4r9hlsPeVUPBMoq++rmBt1ZCpPkmKgwkMKNMNUksnmqsMJx3I/i40x6VVd2x/4wZ
UoN41g0N8IF9Cuky75EWqVe4alLRwvlJBojRSnm0Ij5jaXhrlv+laRq+uNxaLV1IdDaUZoO0dAeQ
HeyTE+dBP29n1U4iNl3KL7ibwjvoOU72KNprLXlV1oRGs5ONY/3RNyIDsswvmhFS6JO2h4Xmz8/0
W4rAQ7m0nx42zB4KtT4FKTVx/k8D5JdkGywt1lz95n21VB/ZXY66CUJjFBqREyRdhOi/m3clNI+C
6FHu9pbg3cQZCOYgyikpY/O7RAB0KMrXGJdddFPYe9pN6uWBA7YIX3qU5ZBtchkdDpfQ6LBnTs2Z
lPtvLYfvb4ERvlkEpO+gCWBQ7z6OjI6fz0hq1HfylpCqMHC+nD9R+Y8C5UCKXx2x5WV6AcEe5/Mu
SuKICGsDserKhLkHMnixzOoW4IpSbakfOF4saWtoHDCj8Ks9dxMyUiU6+ACL/Dm47uwWvZWrLnXZ
fVoqgDkNkXnNR2F0oACanAU5tWRkl7ZftWCPSEu5HSCkkMw4+cT1ErEVnnxu2jeKCq35L9ml+/k6
+yP5XT3Mv1uptMVZkcrXA6rrGnDYoKUHuzC7Y3X20b2pz09b79SfuKE5PuaNV0lnzjOxxhhHKkkK
5xcnEu0lCphlmra8dr3zRIqWAhMSGzlLS/v8JnwzcetOB3ZlYwBkWaHXuTK7w61zuxW+CIvZ5Mo6
zIXcMrbdpRpdwT5dY4T3H1tgCeqOvsphpG6Oa07/+ydrMjOAXpCStEm0AmsUHYuO3ZCs46rXDOS9
65O0u2XzDtK0zOrx8vd0SPY1ovgW7w7tdSTn4Vu02ErUKonGcqFNOvMfH3STUEnsk3LewRNK80aJ
Gx+51Rbp1d88aA4hExdpAQ9wMVpyQGWClumDRnOhbV/jjK98tiPw5ebUfpF7pigwPGh2s1XKMkdA
fsoqfGiVf9rd0bCxT0Amm8sScWza0qQwDWQScWtXWuTcnWQduJaC1GBR3HYEtwriLLh8OMOoorRn
glUSTQRnWrkgS53+aH6eQneOGSUGOvuPM5Nkcjv34i+lDy4jkF1g1H3xDqC8GaOh3mcQRi4CQvuY
O5viijZVGkaHFwX+z0kEqxGlxq09ACfQtN1PAOCAfTaHU4F23xG2wUFo3DUf03zZ8oVRdWeg9w+f
H1P94vlw5BSdE4YgEMKNP5JXs366IWHDTdNmNKEbV9jkFUjui0eERjg2O92gKbUdO1QEq6HtwqmB
1zk0ScYbU0CApkqIueezxTQS4uNaPRg9v5QUjE9ULzBpk/TIpPSeoSdoY54+a0R+/xwdoog3dCkr
oyngtIRpPVN3BvWuwi+wXN1tSxURjEULsQz9WnqN8kBk08B1yqY6/Z+R4yY315bDV/UUDsF9/KkN
eSMZFQcFglNRNluU8RTtyQi4Tx30K7tNkJa15N+klmcwJubAfY9QnOUTv395nunx2jnir5kt01rE
kAFanP9Q5LC6mQZ7CsqMui5FTFamPOyMXLCX37R/xRjhkH3QJ9gxq+hyQM0Y/V9s2kJwSWvffSxP
F94rh4GZ9P7DnQ/EztUAUUPI0BcLBpk//1sDTo0OxEqQ8R8Oan4ycivqpnXycRHCWK/QHjFZnORu
V9AmUGUllhaIF84nKD4FTQHPDT3q6IG5k1q6yhfv1n6f8ahMuZzMNppEJsisxYVVXBy8OE4CwmDZ
dXjLPOk/EHIWA1/dlQqzdMxXy9lh7fAxnBmIMdHZFvXjXKoNeQVeRcQ+Gq82cWF6apMAced+vydW
hDXEWxi+meb/Q8Fp++pYj4CtbbfGquoA1rb0Ryz1d/UEYbW2dA2eNG/C26+4afjcz+RX59NzL1R/
bizAU5F+8d2VGhMyif4ZEMlfFfcFQdRIViVPTTHRjs4IAY4DvAHfUPCduM+e4DQo71BJ4fMv+eta
Ql3hbdNrbgYq8XN5JRORZ14fi4K1Ydk923mdd9JpN8owri4OeP0G8UrHY5w4ujO71Txn6kdAM8BM
fuH25gn7lhFhvDjMN8XwTevhyxm6IQefvomhODHWQyi5oOMXXe7VICnyzzGmGd67GP+HG4U6Zaxc
5GJnrROPwGRWBuyyVelz0C9aQsnwwmqR21FPY5njY/PCNV+WoQ/Myz9hJzxWj0cYmpvFSDpmc3r3
xNxhSeCCAbUkEOdRuami3U99VKOyKiQdLJsyLfV7QDBzsW+LwqgBPNIkb2n8Ep20tSq6TfnnP/zh
W0H/yMkC4TmQ4MjyMd74QDN44k7AEVlkjjaQR/g8a9Ed002rhYNmzNFYr6jkKD6lmHsYXmgaCT3e
E3QfK/S10+6nwkga45pQ5BciW9ZGEKMVlZ7dyZdxt22+Q36UIxliM7nc1bs0bSss8/YFkNLJgfHF
Sjawp2v4luX6H4EVSiP27zGMyCnHGzAj+l/Bks92LB72pCGa3TGlPF1bLOnxfGWByOepMsYnoVoD
9Dn0QVRHe+n1Ujj7vGn9KZcZUuLkT7EYnPjhtFtXl7wdOKM4uLpsqpfA6zZglZBLA7DQrpbwnCuL
mwullOf65UESpg97Od88rcxXy0G7+j+TK42bWzY1ZuOpeqfC8PH0PEM/wQIqpaMIQMzvzqBz/woz
Ips8lKD4otCtBZN4yB8OQ1zGc8PJ3jZz9gH3ZV08RI9hy3jrzu2V42YrNZHS7orRMLZhfJ8to6bK
g07eSXoOqE6UYhsde0ZKIz/7oQ85oDHwwysakvR+oHFpJDoJqi6zRWGG3NYUz8vsLXz/Tm05jIcW
EtMHl1uyEocDnLGjNTYunNDPteWqlWgV8gdNLzm8LUn7VuFQQRV0KGJpGChuxgy9vNA4ZrqClWHU
58ItEWREsArdW7y6IrcbTRYF3mo/+SnuzanNNXKLwk/dYld6APDt/VdeJ0+RzH0Fur3ePFin/+E0
/ZaCAqhOoC34y2mywlRmvrj/kYXlMG4GnjzgkxRYSccm/yTYAzQbDVa5zNpfMc2ft3xoQpoLdkyD
5YGF4Zj8vYl/PmqWy/nuGyI3ffV+QUkbsxnH8PpcUgOWsMi9To4UExVwS21uxu+oiNTdGTspbTM4
xuFiZThijcnynNuGrxPODd8P6mdXMx6izyvFqOYoNB7Pjm4Rgj5aZPadYppFWehAfdx+U8M6gWoP
s7lz9nKvKEsmhgG0SmWn9wgudujXgT7qF5hDSNHU7yRGFRvGnAuSD4rJm63Ln4J/cZzFisz3htUb
l2zkgx1KVPA305BUsI23dSZGBZ7VPzE8YdaCKvvam9qUUIC32u3hLZa5inHK1Wj4423XfUIPvkfg
w9N7uGzCHdWND+4VeP4WCj0KDg9dnzE2UawmfMa3Hjrolw2av2/sJ/VooHeniuWU3nTuoz2I6LpH
y31Pj5oFJ2r91hiMeH5pzMG3bSEiRaLnRCePdiMqlvMab6D4G5TvKnnApaArq8mf32qWEq8ZcMrE
+//1NJr+l7OxgaZDFV6qoJ3tlmIZPUtqeYfU6btnAGifXijNDEaQjyLrOQHR4uPF5KIel3vFb6KI
IYn61wAvBDSk+yP5yVa4sHOpaAimyal2YFsRamdTOD8ryCbdHxmXniWZsFkeBGcXe53REHujEicw
pVFL8lzDvZFZoDoWfGA4Uf4L2o7Ba77RnzxQYNyTWmAulhGSXw1tGJRn87aKY6Y2SbxM+dO94DBs
psphgrLJLCArBoxOUivXdPpOwz53NvRSthnqat1IZLVptaqpxOXp39vUBxmW6S6LBqjOypU7OutK
uD/82jhND8xjlxybZGzI80N5mIH9V3kIfj7ustC1EUcGqStMPTvsgjB1Y76PdyXcpXi1BFd0ugRm
1NhD/JSUAht0vPE6dE5dTk0rcFf+hoXdd1SQKSamZ9lJWzMcXrPxfxGkP7I8tl088py1hTXYtSTN
TWbbL6eCaaDo+rFW8A2IDyQWaN2i1cBUcTYWlJ341ZgHf+Cwxk1vrayORvdYKkQ//gnmnEmOQbKG
Hzd0rUynu3DIXH+CTnv+tHZ2fIBtJy1e+jGXZlwW2BTaetR23npIO+nJW3I6rDA0pgyhSUSQNU2M
y8UMzUtUPxUzVtGniewN/msy8TeoY0IRkmum71gOL9RkcbjuXmiHLgnj/dVO0/ZNkCyFpvrUbmdG
5zy5IrMjmYJKNLzx4uMywc70yi4ioDGCR39YLSSz+CwN8k22nQoyQd8VOxuBbE/86IBIkRF57fKF
h9rnXM4GiDIRfSSUnM3MO/j42o+vixmNhVDwsydRrr0FqSFdo3oWSutwtn2P1+bQem7rD9BTveQU
gzFk8OS+nVSZeE0WB2mkBNfVNNT44giygmKZNdO3HSVQEy4INpQoni9DWNzPpSV7WWWwefD6vdsS
dN2wgbEKTNoriKhl0CXMNi3sl9FuwaWHFp/xzoNvRq91VM1C0I0kJzkJEqn5QPDkeb2ZE32poim2
xEeXpa2gDLK/HJ3KLxMrOOWQSVWdH7iBTJuqbZnOhv6eWyPt0F4jdv014D+PuI6z9niBLdjVFYA0
m3Bz0bnoAtABYUFkBuN/CRiGglMM5YfAQC2e5RClPPACKlSqECWvyaOnpO6QkyF2Zq9C0D6DCDdE
OAve0kfN/HrY27hpSU6yUBbSZFs+9Q3KBe3tCtCSBN1YRgos05AMyistg7JiFNV7ub4FwC3fD51K
Q5TOKA/n4X0K55tEc+y4fyn31Z01yrGCwfU7llwcrJdkhg3STfPEqupw/89jhiUzahbvURFmtyni
N4CTUHvEgHrPsSWUhDsscwfCAeFSGBRqL6crSrKq5z1hKYE2b2o0g5IQYkh3YeZLEXZQutFfMQK4
a+jFgSbcHmj7jZ5techR9UNgmBb6ICVMdEe4Byqgz42f02hcw9XRTLNWnbx8wZQwnD63yPOF4m0Z
Ph8svstdXAhT7pVhHc6FUgNbGXzfq8mrSduRideTvzXDp6mWlz8I/ccIHgujo6wA/GRPixp+Izr4
o/RMVqdAc+WQTcnHiw/xih6NKiy2nIfz/kDUi79wWuBiMd2MgilrS4ko69Hudgzn6s4sW1cyqqH6
/MHoSdB7OrcA2FmdoepLxC1rL6qaux9O+/8FuDnHGFqz0yz67OuZJxmnQgiSe0hiTiQJAXZFZeC2
JQzD1LNJvf0wMSpr6SVoHuY2rByhUY0TH7lfwy0gKfU4NS643KGhB9unIsqoeoevcPdSwnvKmMbE
/T5vzsuDJxTuotG/N0ArbvnDJfEATM858p1/7TcYdhJGwk73kAGxWat3ydkqMqLdXYTL2RklwWMl
wRy5Q17mKoRzhJzb+PGbg8HZQbivD1syvtNSpj720roB4fFQ6S/+zATA1R+JYv8o2b0XYPt8DsJp
9muwP4A7iNKZsnsIupmyMmiLqIDIZHtxi1Upss+JVHO9uQYBh5gqghhDOoW2kL/NgBS5klABN5rp
groH5H9kXNKhWLEXxpP+UdUskz2J52Zmj3nbVP+XRD6Dnf+4UnIjsMx7zDORwXLcf0ye2piBnCOx
7S4jQBfiR17AGE28Y2deun4c8BzZp5iNQacID5JLjsX5uqBusSnPJ2N0tdR3Nc9Ts+2VYx3+NtWp
HIxW7Vd/E4ndDM2ZKTI8NA+1nwiNo0gk8SpiyLLDpekTz+9rhIkdztpfoLmSzZ3l8iB5bOKx2X5X
ONFwrEUhsBFLaNkgXTKe+7uUh0j7sxmxtTcj8HYB4XnBTpXPr8FnqRViK91c67Qg727IDdtZNTlM
LIwABGB1U+Ypk5JfJT/qML12LeIGLsIwB6ut7W75Fts178jJNsJv9m4JEWhWy7DqjXWpLal1fgx5
UJnSlPVHR3rtVoFtkqxF1f3RnsptMW2F1oZA63EAIODu1GM+wCDgOqACl/Qx6QAmI+lssNjwP6Ox
HXrXlOuq0JysDizZERFbhRZJhPxC/DaFMIL2GUydMGpfdUxrnSSJy4Wx6BmAQLWflZNinFcV/pQC
K6qCGhRbDQ9AckkCivkRJLPttYSslWo102UHK9JXPHdGRRixFLt9i1S12vyOvugT8YPrv0iDFbG7
yCSYhhj2MFcbwqOjdNWnClhR8AS7JP87J4TodDuYVqOW3garXcsxPnom0EsvGjFtovkzVLhcxhvK
UMMOI++Exrq+i3uMf8h5lFjcLDU3Fwq7p/QCTAvXGu6yKsI3kllvImO4xh4Vx4R4lIiJoThHSLbD
YM2YLyAhwZ0bhxwJRs06lTQZAk8ItMU6kBoEgfCBnxnpxCk5G4QHh5WlW1U6QstrxKaZpi7BjSTa
JcLREZLU+h7EEFd4gHm04c45J6OiRISZMckzLpk7UqMaj9IRJadD1NSPH6+dKGJ7fXuTINBWjxZX
qEbK1Rwx2xYau8BbT5r+XbyKtmJbzyaiDOcDlYHBS6bqP9YGrQaWwooxr5vDAToEE8cZYa94MpPw
jJoBC5iHlPL5q5jwGrpySPWt+0LG/k5NGY/ZhQPqchO+c7vKxwRm6fLQ5gicTNATSvHB2WmDjym0
ZDI481Q8GCKA9w+VpsIdvyyD6VTs49dfVldEqmhJlvUdf9ZXHZvFp92FugDPjfEjuX6RGKHzcyh5
AWAccS4y0UAnHvWJRXcJt5F+QArqGN8SaNhUcbRmRDyn2QAddx9gSbkr9tM/d0mdb5sCjrUHXHG7
LK8XlwSQLN/H+maL1skZRD8n5mNr1WCejQ55uRefH4+aLIZ0V7a8EUtD58Tw8sd4PVpS5vgX6XAn
bla4pAYAdwkb5DVyQEeY4y3lfrXhaKjTKehe0oXI06NGFS0goy0gsQBpYWrinGQuzs+XoFPE8oiS
f/PyLTXcFbGnOPSiYRSge4OKBJcRngrW+egSgqdPbIe42v1/UG6t83mleMQcD+0OW0+KFicBSm7H
XZXLVOr99uvwKSnMd2NsY7PS5yiE/xwcISx3SMcdDvgIyuGtIw30Bk4CsDFKkVQ3xjtj7vd6MVOE
/Wit1ZFV5qZT5FimUZ+JVR+GMe9PoHAHEua+BvHZxRZvA0b7G9QVjeBz1YupMt/8XSse4LS+jB3/
GS/G3RzY0GYgTOIY/apQzF3OU8gDq1CSKONY86YSW//eIFwB/aSMHMFNHMJszti63BrUaW5gqI6Z
V7221KR2gHmB9jRitfuUlp+jAUtAwF2uT2Iu4YcnhBIvxlbS1uY2szwAxNzqhBAV3juECEO9LksF
JNYODXNqn2gg3ER8zGOwsLdxJs2SxfhcdZcn8JQ4Z2BE47RbcA8bwjWyi+di6ibwBhhYY2lvyfyI
qCVVwtwZnKs6LoNJG6R55kEf6hbbTETj0mFU29l1OxWg/NylLQIDuhRdPd0heo/qQEvrTIWQi0ev
61NUE0q7nEdfpn4OZQIdCu9ZYrFbn7nCsGyyqSDaB7KKsOlnMLLiRBNG3Ryq4xByoYNybHUcwI+p
Y9CqhQo3YTbT1KTWDl9/PTKXZ0ll0A6p9EYCWWpPwRDvwHqMUa+QocRiLkBkd5/cmp75umeTowTe
WZcNhS3OPJ2B6hFgUKOlk+jmw8akgx+SM8vs+hxraQ8fUVIU8T08RQgjZrsNRMn7VheSRWLctFjh
NE0TP6k6oJtV1uWZ8VJt+86f1hRONgjoPSHXVLo2sZnMPAqh7eBs9nYY0/MTfseTiC4Vg9mapjca
v0NaQHWZ1TM5z1mFWPvBtH4bvuxTa8xwmWDgBVmj3GNBulkNW2qvnao2b6Q02QO/eNAe6D9CtXFj
p+YZJkhPz/XTXsiTT/LKPyeeq8cI8YtIy9VJs92kZ4MKx4uHe9sekq3nEv1T6A45CksI2roGKhGI
W6nnxXA0+LsM2sEo7kRCoFO2n1X9xmeJTl7lyN4CHTSr1sFT53rkv6GbIA1Eb5o75Bb8atZCixNG
4CHSL1DdfaiIYvUsRs0NFsaCvC6xePa6ZG0+XuJFzXm9bs+UKCGvbCDsTdSni2B+LKQ3DanPocDZ
2Nh8BcVNpcQGzk0korEBDPQpeMUDC7LGbIoQHVnsjb/cTdY4xyGGqHBDpdLlXbHtMa94VE2YnyiU
lWOa86/nZ9jbRyuNNMYScSmyAm/wtuhhfKWA9I7mHkYi48K9veY2eYxT7NeMX5EwELhQ0U4nStAY
kKQ+Mgsz57FQMUzjhL438JhFLmwHAhRT+BD8adSNTyCfzsqD7T3sCIeRg80t4TTgPOwB0Cugx3ug
uj3kvBqo4rWnoE3NuO0ZDuGICi41VVaHHhCzcbZsPHXQGip9yCW99bGbpjecETACJGCbTHFuI0+1
0tF800vC2YCjBcN5V22MeDVzyzhxHaZEoWyDs6gCMhNv8FLgMOccdnQz2k6fbmF3XeNAK9xw4ju+
8D8rFPWAZXPJHDhOjSMT3otrSFGh7oi7cf3Pgx3psKBKv8AEgClOcZrpZR+RVP2SRQgtur+B9+6L
MRBVbrk8GfVJrCedfuBM15FKxrYQIGA6EC+y8Zfp60XbQ0jTd5p7vnYYfKzK/1Lvg7pLy7c+h+r8
HoMDr3AVWbZr/4N9e5lT36HgfdKcDre3SgbHLA7Huur82JHKjIdO4yAghshngpxGWrBi9c+5CJDZ
6Zm7qHypw7EcOziZ3TlEckD5ZzT4DEoFQOU5OAUruvcULMG1j69+M3ZGmFT4ZIwF5+qrr6M0bQ+o
vKn5YFmuyZBxVyCkbCchz2cmMPqQ3+V//C+XWh+lK7yk6A4UyyZJAOy3flFitQanoSTVXk93CgN2
Mv+EvJAtfOPJDzb6WeeZEdrXEmri4A9a39JEhfFFUjVMlnBwY5M5/yXZC/reBduqw0/3o9kmmOst
+7WGHu/5uL1Usd/yKpDMokLFxmQcsPYjpTLnaznDsODAHz//E8fALOWAvUNJLFBYXVnMgswl43sA
xPYlZMGgfHqZqlpeAA/aBfe3voxSMxSCiq/XryjpvjZkLwuBJBSLQN/F9YTh16g4fdfEdBL0itkT
HErWBl60zBt91wf9zMiTeWbW+2AdYs5Yhl88Irw8T6usFOZ9Mx4u1VYiy7EyBmm3GseMbwMW4EDI
BSwIySDhEcI/eNr6JMlWgTpM3nAVhlROFqghbT9ZAnrem/TZyoCjVTgRnbB/JY4yIaaACQQ+27m3
nRc9LghFdP8dbYaZRndyMn6TxcKOyFmC/ytvQf9al3D66B0xJxrkBy6bWvbHgFQOp2aqvLut64nO
3bVNdqpX+cMqaeWaEdu/LJGP8Dba/urjvgbhPBXHx0ErSYjQYLECOag/5HnKeSSI6I0/KsgDzkzy
3SMHHZcAXflO2Yum2jTtvoMFvr8mvIGwTaLWe5417j6T6a2bBPcB2cMy7vZqw/13FQ2MyVCzyaFq
YhjcrDNEsQgDLxPpS3HoEfP5xE++hBAvYT7/Xj3TZTgEVuMyduJdmZv9Lpb94yLG8U4XjsgZvowR
WFEbmi99LW628EQ17WeLd4REa5Y7+jUqtAjYdSP9Z9DFLovt1R7Zc1/v1+e1B6TJEHoxcPr2bxMS
Ks/CxiknMhTzboJX88WRBiLuIXzPhtan7SshNj3zbDZZtTmUkudNC2xmEno3lCEAaEor/UJGXIqO
QwRd0B+9Li/SOK1e+O9tLt76fPXQDSV9TjfVUo3sSpE+WsH6bT6yfkfQZmW0gtt3fkBcWlhXjIWq
D5zqgtaBJkR/lnQL5eG71kTE/coKF+waFY2k4Hv8jNT7GI9iESw3eg3x8lO0uETzH6HxTN33VQZN
Y42+C24Z18eCJtUHhEIPPaLd0JoX62BwFQ8XsJagNd+nvH+Oxd9PARgE75teDWm2oGLA8LP2NpYQ
lvNVMNIoxpsEiFlNUcKsxrAyioe+3cd7/1ASjL+ToKZQuwsevl0ugpQNTW9S7MuYkm/y8a1bXSTz
vOrBEQDZjGyBeo1/q5uo4EyNCRMJ8tjZZs3stzKYGz4A8RFnfx9VvXwNSBPXmTKEqiRZiQJQVDBl
EjtDSkgqAFTZhUWYY41et+4l7UkkNQp+Yu67Xs0O2fL8TO9vE6Whhhz+5ZdMJSW1KVrxnePucmC3
kFU7qGgUfCT2Nwi0uQmoLwpLECumehK8K9n/QD/lv8HZTaGmtXiMnmkRBiYyWttxnw8f4y/gGutV
aEAlQQVce3SBK4IHH0Fhw2Qi7XQNkbkdOJVIiM0gJxulWt57RhTZj2p/5TLcTVoQ9hLzDlw5o88o
kX+otL28F+gQZdcZA2J1GOI+HEk9IT94xdO9JIEKXWDSf2lDvElEyjVUJyA2wOvanLu8JiHslSsa
WlCqhDnATVK26nzlfCvO17SZC1sAItagI2AyhLpfLlUi7HyeihmaEImjht2C/5B+7nQ5wr9Clp+U
KrW3Xd+m6KQ14yQhbkIfq/9ms6Bdx5K9M4N+eAvJEhwEOzwwefvR+pz/LzRCjZHGAO+UmmXdCL66
bKyxsnYYjflp60mxDFmWaft+NTTepCN3ncvWybyriMBqdu+HVMqZWYTvevD30ihs8H084Z1fz82F
ZdDAqdhNyF/PToaKxPrBKMK9r8wLiOdjjfWRYuYPZoMw+vpuXNM1L1off0NZ9RaBDyvgA/esSdY2
YEhiithvWDMrDqmqc8er5E+QEviO3jcNu7kdSojvaQbNCp1mHlSrQkuvHZfHbVTWq9EC6ceBUEZW
lE0jvdSka/3gRZWxOXQthQhMF+MEsZHpRDJTed5QsxANFTSpyPUKF1soj6Mb3MLQI618PQzEq2ZC
gNgaDFHbdt7eglTv+GIRdFUD5iY3764pfU/WV+GqBLzQQxLNtyRHIfh+l75P2W8jRj4Q17IZ66ou
DG7W//9R0uzgQ8LMfccN/kXSpqY1C8HBkt22mN4yEyngaYrO90bHjdQ6oaW0bEFGhflvVOVp0GYm
8QWIjX+wfSGm5BhqVYadvnEiyzzEQSOC42VvlrIGkrDJZpB8LiPX7hMbfQjGpMIalBeHr5fi8P/B
PR8tm36t3z/E4v6AcLr1YgKUX+tg4oDklZt7zxl1/vUZHT2t0Z77owHDii2uJTT7G0ZwjjrLR57R
hINioXlay3c5EEAfoAeGD03twlb1SajFum1L3YeDV7Pi3m3na7UwqYoMGRSMEU8/Ttl6FngY6upx
F5v88Q143A32iNfdbNDKvvmANcbNayC2BByOIos5onzZYvbRbxQOSOyUBlUyQxEAfbI0t08QqaYa
8xRFf7Vua14/Q3UiFOc704S3o32GblSJ3A+XoJYedDRdkFC+VTz1Mj0dNSzC5j8h6UB6daT1mf1E
Z/j9iOQc6Cd7RG6B37BwNOZWsPvyRPSrgWjSKkWSv6StSquG05uCL4EftDDiC77/IDAE/Oik2R30
AyVDRMgm3kL+eEKkJpdeQwoSUOlc1cxKGouSfW0txCsCxGPDUwolY6JMmGNlXfmeSytqPYmfQP+l
0vXh0Gs6yPZO2vq6oOFH4FimUEo7+I2uufDLAvKEGtJWSun0MTQKrMgLpihNXuifR4G3Jtk5IxTx
Q7pZiR11T2WiCiPRl49iSPb1GrcdjkUwkuGJvy5epO752jesQRO/GxzWbVuivybxz8vO/WhP/UP2
LeS5qF9al/HGYZZIHI/J/85xtxhN1VpBDeLPoHusWHZwLbJv5TQQSlMcuKbgxuPJ9MXyZ3BBLnNv
9jF3MMuuTaQOwWddovfpikngWHlq4qr7ZiUqU6uXGpZcA2UicI12IRTnNjDPc9l/a/GJGFKOb51z
GAHNDM6r+s6UVM4Mn1PT0Y19mTkZWKql+1Jnpf+lvd7e/uXYV0MZ5xSHRAxwzOSzUM8WHCU49Ssg
ugou8Vy+omk8ZQRYL59dKFLkDqexD5zoSmCBd8PUWqzy27slM35swk9pSxy7xcWiRnxV6upFa6/Z
K+FQElB+B8zME8e3CBI1bZ1rf6aZ+Foea4jt4o4Jw2qznPTlZpJTVbyzh9t81jq+bNMKuBPCZKCo
9q/2QzbjZhlxX+PQmV8EdC+gN5Ci+zdIXT7vUKRWwN89jjlV4lr9bD267/IFoHBn1C7gqK2/r9dU
L3psyK2TJRg96kuThwGc9TSFAifYK8BFMGAF/nfdIqMmbB5R0mDgWXAPjpLfB2GXh9JaRflZbw+B
/epLXd6MP5P38NUNG+3SvsPtdn+sGDCBKyjFf9du/EU46LvmN04uPg26pfCpMT0iotgLjIqODn7e
m4UnGA2no8RlLqela3jPidjie+ftLMbKwmR8l+wwAsZFsgQ+95pP7H6EqIzbTcN4uRD7kMWeQNR6
AfM5LKDaPqspn9NURyEuN+gUFauRzEo/XXzGCwwi12qZ4HSa3i2G0NBwYaANuS8CK3r2WHpRZc5B
8WByqJr7BmO79EeStlTUedymTlKoVuNXuts/fyfb68gZSHYJNu4JnHCy/4gQLkODOVm45CWyT3Ce
PWCjtnasSSntMO/uEm52sg9O2k8EBxY/RpwIiL/CcD0uWtFZySWD1BcHJ5r47ZE42YN1LnenIEwS
Ym9v23IzflXokjUV8TsD+h0adk8kuv44K8x5bytH2fEfiz8UgGlrGHh8Sak5+sIe/BEr0NlgFNJa
PzpuioUqjcrzLq+gkdrne1Uf6M2JTCGXZs2eOhwlLYYStrr+rLRMtHgpW5yTIKYhqF5OOzrodWMu
FQI2qXGsDAHYUL3MWbmHBI0bG5TKX84srH2w7twe5pjXYX7FvcXxTSiXqYZ095rHIMNHYrsHucog
wl4MxqNkQiEXXIoUWLCs9mnYyKX+zmphq31+IvtgdmaZAK2fNdpbvLncSiIo54oAcL8uLzSn92AY
oQRmPP7Vp55eDMyq1Md6dTAwZ2R+tSD+vq5zQlHzXX1KwcMppSJGe0SSHLX8VVGXvs4ZKVSRpjr+
IjxLkan4+N34ssMwl+5t1qa+z20+LtBo+dX0VItZevbI9BQilFZK2RBqjMlPwcdU06O+An1A3cNO
m85gdbwe9zcOsNkhFBrw0QhHTnwtWIMtxNPGx0B6phXjbEVCkzJnBnaDV/5nvexsp1xWNsDoZvpo
maSNl22mIDO2mT1t1XFm69gr7UFVxc0IOMIjcafu7o4DGAwS4k4Odguy+Cfk7jY3BVlLIHuzo72z
oO7/Gt4NcN8ws/PyfP8+DQsghaFOdUvkn3DGwYdGM6hUFHppgoxmxi/Tfqnrlu+D0nyDWTnyHNXF
Ha5SgvmdF8vm9wMM9Ql0QOJY83kOy7WFn6GK3i0wvEZEQLAjkPvhSY2WqLA3dXNMV5PEfhSpnK0Z
gcr+1ZuhzgdM6DuprcWTyYA1nWHou62eOokX+6a8SUuriOmPEBZACLhxp+5LPPov4OrfFef9VfL6
JzmyqyyYUDkzKV8Kfi+cma6Fkybt2bpWF4gS8ykNwoEnLDLzpC5HdB4olTA2buZJlIYcKmwUzDno
tc3IxmgpiI2ZhM34aLls5AX4ThEeCTccHosd0kg77zW83vOT7Wcw9i/IOQa8i66UqBgpg7T9mdxs
1nVpT5J222qV+SC0oJ/HTuG2IlB+a0ZU0hVXO0wl3o5kg/cPmEFNLNmtE0NOp40Xo8yHdXaqB8if
Zxm01NkXbSdMR0PED/7d/9EQe4NTd06BHqkDFRfGRwhNDGWGnRp6zRZpzrAGcdXCEdO0nkvhb4Qq
2p+OvgABhztqlymJlu0VAKTuSgCls6qadAxTRGEnafVoyMomThBIviNLMH2XYPeDzMTCR4/sbFoQ
1dzjagZzAle7fUGGOhoANHoA9ox3/FJU6boUNB+G7F1Go556ArbuswTHL72l/fXu7MT/iz0WvEAg
BhwxMGnLHbLx/RFjJRBEoI4FaiAc+xJuSowGSbStZu9wvGzbNTW/WS80kmP8PibsSaQtX6aGyWUo
+uGpRE+aWUbtwcXNv26i4IFuephVekmB2MAMS4ktCwPRF5i5IUfsGvVZe4JpU8NqI0JSiGgbzn6m
RqAy8mTKLhTRUuqpNo98QF+2g6r2D5KCuaNEjT+P8FA0l6qEVl+1P7DEkf+54tm/R82oi1VNKanI
AEj+iMJwiigRHOCHHSz/67hiezW4DQd669itdRERjBPopq/ATEDUe/NY06DB9bwm/JFT+C1uj8nR
3HwHBCcOK1TZfHCXaLNyqEe87Xo3eg0ZAUDsyzVsv5nTm+nXcZyBzrJ0hoqlOgYe2joQCno7fdmr
F2O4I5JkxLMPakNKfEO8w64jnQpvMMc3zDx3KxQ5rP6S1//1jpLfF01FIBvFIrr3SYu69JD9h91t
AL3ybs6oZ3YrStlSeqW/XQug5syVi07Iov4lyPROtzhNbnTaq3JmfVwMDwmDyuS8iOtJhrBrJKf2
ZJKDYCEPt+Gmc5ykLUj4fpTfx96LwEst+YX5AvDvhj3L/k8ARHEIUGeN68thqPFUQ6T9rzNpuKVo
xbbYUFeY4ur4HbdVouJT3dYEDX6URVwTjSOi1WaILUHpuu2fIpq62mEyOO4TGxvBkYOhZ8hx5H5V
s4cyNX+Hm4Pw+Wq9fcAVef46nUGKm5pQerqiQYQMxKfxIZhmfNL17VA0kLumz8uDBeS6IG8BHlL7
P076jiTjnS8qYQbbSD+QsO/muRlaVj15zX2bH28oRjg/Ftt3V09eEBgSjwpk1z9vMaQpxobod+PZ
unSs3lmtCxhxl8fEc7CZIsSJz5wYwKeWqZZpZn+hdCPCoio+KPJCZE5nvguTHdWpx6TjurH4rpIE
UWyjL3c3o7TvDNGo0byjOmhwjU86cwa7QPi+0y0T3WMUPFQhHBJkZOIzMs9sbsgNqSHFWOAFQokZ
LrIrmbQT4FJQzuMOkXXFkxcy2DUiV4qCwCzGhnfWcIN2ZGIFiduDI+rpQaX0CSOPTo0dK2MEQMWy
mqbLSIfgE2r/K7terYg3Jjk4q7tyjSLlAC8DUr0HBbsyXkHVPisQkBhjw/FZrArUdKGu4NSnb3JZ
wUir5sc+mww/3ieTc+rR9a/RzRh/TWWkOHq3v25OHbuAynixVl1g+w1sF9tDjmFXr2qw+hTzzms4
mhBXmRuICnUq4udbyH1adHmH61j7Fn9EVe+vp3qeVsHDs5zI2JA0q0zZTDDEWvVvxOP5PUvNBPLa
CrS0DZ6DiRX9fFvIVxUdlm4v/ZJk2xqA4Kh9CXJi+CqVb36y9WNIXUJ0uHjNNUF4pPJxkn4dL8SF
GMTkvJf8QXT0NA10s0Q/4EiyfE0QVVh5osYvgpAJ1UC9OEG7GiabsG4nPA+RUHN+imrUeJUS6DzW
gaAtrrykC0QShvs3fVw2IoQrTr6XPWey+MMpJ5KePGSdxXbOiWPM2j6svYNDTzvbY0m+R1fldX9j
8VNT0ZGwJulGkfaTS8p5SRrMFLj4XZh2tDfJxrAlGMg6Cuf0l8NSKfbcWZfqZmPSXBL76DttPXe2
x2aFhGgRo8SRgG5O1gEGYuSeP5wPttNAGpr9gtSw8qAOl1criOXdgZOk8EourFUsutgwReZH/pVz
lumX3mKnFezAN2ASmzhQM2hjboe9SbwijffJk6i7ZmGnlJGp9Z5Yg8HBBlmvuFE8S7T6gKIJh7GC
tvNSRpFpbKEp7UyTLmREDk2s8rsXScTwj/Hbn5F53Zgx28Cr2RthjzYcHSVKbPGy7ahU3B0Xa0tW
cyDvyL1r+xLjEyPsnWjo37mQeCbY1yeYhZzI0xKxsRXnCcBcIMC178xRkoyuqRjq9vtSwMm5muYN
fVLhiKzQaXgDkKNakGqX6a5QbxvQLdR/SOU0Aq7ACgUF+5SqHMsup5WLLsKXhEZ2s8Do/pcci+uW
Yc93a+B68g9ZT3VL4aCg1WKsOfHE9e0CmmpWRE20OdaSZkgVKfdHs2iuoxZU5egWjT//0IXjy871
dG6ZBNHjkSGaZkBQK8pqCn0UzTtPqPoNwT5GSKREc0CylrN7B/YrO5JNiAtUkzWOppjPnpeb4RDs
uEThNQQDqrQHic4a8Xsdf85DuJkptfmLfcoxac3BHlbUbuWVBzl06OzAyNM2qRERPiYUTz8stmr7
Iv5ZM4LmFWbfc0RKeAiysKUhAYaTDOOCPDRvOxRp2CQYTHQKgSPrJxna8HFQ2FgCIISs9zyfiHyF
OFG+1zMr1ecvUU5HnUAY0UV2FAACkC+Rn5uGe48rfX6y4iS7kjZsF8rpQ/+3Tvm1T2/Zy/+1Toa/
HHoRfdo7OA26cMVV8NCoxO1J6EiWe2yjR9PqS/NBiHfOhvsgnJByTiJWDJKGBvESUrEi13us4nrm
9sZXcr80T0ATxzxb8r8WEI4d7o+rIHAW2iThd6zU0S65Fn7pVoVJKKi0p00xl0h/uoQvcEyMWgoe
Hx63cOLI5bdGyGANLFs8i4nxqTwJuRxKHbfm7+8Kvgu/VB/PSwZrbJOoX9Y/GGiiWq3l41aeOrKM
MayNYeZSO8FQKEIVyyNrd5gnoo5E3oGc4NHZPH2bKkZIBO2Gdd1IuN2w9dPaJdmdpuJRg8nV7QZA
QswGrEHRVsYRSbJJ/jV5CZBvEFdY4LQuhwX0ommYGHNlwy+HEZsuLfrDsz+CLISUSaO3jjI3xDKS
PEC84Pk+LlvAFmcInM6j1W0HkXr9ZzRlcDpbneFeW2jl0r1LEtfCJ/wdvsDchhvKff+l6VPyDjlL
6OcNn/ihOZS2mPqtB6rLr4sR4B0q1sfD477sjDI5Qv3EdUuxF/lmS9cHcSlqbh4utBfC5Ja5yThq
vhQI78yUORe3aSazaw9JOmT3i7kjnWij7dr3Vu5EtHyFWXtv3cqRHKfWRQ77LUi/IyxamAkLP5ye
N7IqV+odWBBY7X5Ptrav+if6n+lnAZsq0tBtSYd1r3AmhqrH7gztRo1nBn57VEyjLeXmu1MVMgvQ
/W2W9GJ2R8hNRuKx+1rakQQ4waVXl+fwT4izm1zKaw66/KkgDCXaLQwhlycrQMplbI5SnVirrlso
zcA11gY6fJxEyHx6RTs+fuXvWF1/BDLDULhwiE+6nVEqTUZGYTkclGH0FsSQwbLNOmPPKiFQmP4h
RwyKoovXDeEMpbSOK1Atp3LJkkvIhivrsJEk3Lrp91yYaPHrCGCK40KaRS/QcbjMTUxx+daRvHW8
NvU354y1Sb64fiAM/D/uwKvbAE4+PnY8Op2L+i12qkVK3TKKBMfxJdwzHxVq6lXCO0hksTB7FyhU
N66cY82zCe8awyRlYnhLboYcsPI78TgPSQfDu2Y0qqxSgCxZnZaGv0bWko92qmN1//9dyxyzcppn
tKF5fnRxM1J/HKkDO/4eNcO1hNVuS0JdeJo4Yj4ikXigjefx8qguv3O6jGfBzYO6WAiiKLbPUYk5
oi03B+K6hZBUQ6hnDHXSUGGpoI7S5aVqljlq73PAe+vGhT4BCrvcNEYqLSYBARuqcNSA/3Qq33a+
0F4MrKdxpAGY7vWPBLfY6gMIjybXgEZhA1R5QmQtlJufo8RmNACu9VX6AuYJSDtVc1c4zwVoq8Bq
pvN7htU08hLPvJUZPG5SsanFAwxeaXQkpLq24kKcc4NSKT44TTHXguj2QlSuA2M2FSh3GYoeyX8M
VwcA2ceexsAlnrtCntKS62fy2AFxoUxGgE9lvmMbuq8THwYFRazoItNBjypkcuvEMiXNPZWKIu8k
Z4Zdaur2SWbgRdqUGJ9YmBSI2CpddA5+sqKE6HQD8x+aPyFyXZ6QfbAaieKmR5ao2hOp/lZr3zu5
GdTFW2JZe8aT3Mko+QDfGtp1yJF1C7Qt10D63Zz8T3N3O/CZW4GnxILmGq90qRMilk4OhVgSWDUc
V1ffe0jnnM4Y0Xqen7eSFcYzBfRxLFhYLGS52/niAo5owHBIlp1oIqRQkdIYqAey4WGwcctvMyF6
T9NA4zNoLIDadPQ1XtWMv0je7OdvtAoXEpnxjt2FtbORmU4maXPIsJpiPhKEnjhcTxqWv8qWF6J6
m0Giur0szBUHgxtzKhjveIvZUIYqPx2SwvHEpsG82pmCGCh8UkbkgknDKtKicikKNLRQ3Z0XnxXz
4JQp/i4V20dlKOXq7/n9iOKxnrPxABtye20ylawUbCyhL7v1g405E77erlNGQj1MIM3LSHYqP9Dz
knNZnvD/8LsxBOITHeiJAlF808X39zhb7+v09msbF0WJSX4i2JEnZ3mXf5FYnljp7oDvcqKnE3MR
FccYdsR0feAfCEk5EK304yTLpKSFPiqvi3mGcgtF7spobsZIO30SjzF+XgCZpdD4l0rCoVamq/Yv
HzT8tZuPk9yyKpqniOljz9yWcivPIzDmk6U4iXX6q9Gj9+mE1Mincjqg64SgoTop/EzHORFX8FlY
CQ6UPBlSQcDcGhCsBKPT+igWrmaHJF55NYCnCQQpNTRs+piOk+JCJSAOnLMeVOnPjxEEIfhjQQiQ
0V5rVHrjYmxfL/Edk7ZJcQt+uWgNevTQ8Ftxs5237WWq5NSl9fWh+eSWefh/YR3WizUlhpLD2AoC
VQIxLOYJYPKoc8RFUuchfI1k8pR2IjPlSKAwDT1yWne56KxUlPCGfnXwsBNibsMLux5qVtnPOHsb
FEpCdRJnmIB4SP48YEWzXHugBi53ogMgaa/goQIs4HzkWtDxdqoEm91dL8bCdlwiiS4VpLTvrOUn
k+UsPyvEXWKIe0RquIk8oL/LnVs/eCf7Yc/j3fKY4U8pNJcWITtMKcRjRQRHI2l9Z9ztzaIuqL4h
y4vjiy/xQWEM361vdR1XaCFsksd1ane6UXuRebBTgeGJGBULVTIqlFCECcj3uwwPO8RwOEUt7ia5
A0v+sPp/1K0M8P0ffzuo+Qcmyme/Lb1F/cTORO7OvnsgN3qTC6Lfj204K9hexguB6xGJUzhekUvW
bqp+zcNDhhBuzWx0wUDuT40EPBolyGDmknFWBHe4b/QGuHXdcJ1sPaP1idz/ZyFdcx89G3C06WRs
pqGKoelDMFOPtc4jHIPZ6n4c+jHQIrUik6NLBnSATo4rftXoscdWyf8QbOGYBssOEVBU+4LqWrHQ
6Ujypr/mLFGLzS7KJ3nrf03k+UQFLmwrrB+1K4vanR0+GbX/rCCVpu6evDExSDxtHCtYBQhpQ6Sw
l+muzN4O8Z/Dl3CZio8g3vXheiEvfurw36OCdmu6rg4cUYwtUWGEfAxNeNEKGO9zl4+ngPqVdssO
3sJ/4yeKOcmLuWiCB5O0cF/nSngkEhdSPkWHMqI1V8W7G/F717OfEzpIGUZOrl7a3xJ1KDcpxAM/
n59jPKNkZJzi41xKs21ow4GUoDg8QF0wI1+FZzv9McicUhQj3D64D5gZ8XRoOPE0oTKBpD5EO/DG
lnLM2xHL/vEAgD26m1A2YRsNBEe2LRjXbv+9ubZyPFkaQV1s0+o0lWkfW+mktGKRgwGOEmw+ux84
IX6+UDWwUt232zS3nTLXwhK5Jzk1/+mSktQ74H3ul2JRfdFL0rGhxo83THgiDROnm/1/DvG3cw+A
Y4L/WIj0rt+YEz8o+dmFT8w6aKeraHxKsBB4Xh4YpKWKH0CiocYr2NbzrUYa9JTuC7ngE3wdrzy/
yyqlwyiGlIvf2v+H06Adc3YThERX2Q3BAzYMfZ/+Ruz1Rvu5g1Gt8B8cXdJA74swZ2wzK5gLTEtY
FSY+5M6Zkn+HSfGUdW8AmBbtB93UBJP+SyIs8IeKjgUk5lQU2TVZagbqyD8liGb1ZMzI9oxirwbt
UNl9HXEt8bNsnwUFoSz7usbIwJ9inCqWeXc4yA5JZCtI1bumINvy+B4zMQK4OREWXe/dB4W54GjI
aCDNm4ueieFJVdsQrc32JnFFmv2AEj3lk4OOVgv4QT3ugCNp93etD9/hZXgr7y5u4E0m8CQRk5Kb
irTYGfN5Xxm4Fg/LGCUt4djr10OJ9U+IrGZUvjONavrv1zf+KkFw8+Mtkswnv1h60bJ37UDq8bA6
ik8pGtuAkQoKrYfnNFvYWZ+DhnG/xB32YjpoB1i+DVqybf/HNr83tbFWvkWsiv4wQZAnluZpTqCc
lgyw3+Y2OYNpl6IS9BPZZvR5WsVvU/yMuTXu+5qCp5ejk14ZieM/55ru8kB2HFYy9vUx8J1ysttp
MgqJiYqU/4Zky9a5vXzBsRHNv0H9zvUMUGuyGGHcy6lcvG2OOpwY5O8dkCWU1o+2LcKlajrFUEtD
MoOMei926UCFlIAhmAQFI1lx61qRgMkYU8fEuzeFgd+BWfeXr7uPJcB0Y+6oRKuBhm2b2jjnpI6S
YO/ZJK8V6v8nfR7XAzmq7gW35FTpOqGKMQ/mAbaEgEObnUrjM/GJ4Oazt4lr1mVrn5jyS1431njk
GX8t0XIWSLlAu/XGGYrmvZP6V0A/A/+ExFDP8odmu4UrITTJxXei/ac2ZwinSAE7sxYsw/KdARVM
CaNPJwlowWby+QOq4wEHJ6XP6BxogsRLDsQgtPo87Bv4/oBKRsHJsD4Z1xozC3dI9CWvLz8gxdHl
2u99Y/gocUKmqkHhQ4tKos5cjw+dRqEppckR9IxI/Ix+HvtpzQ8gxqCqAh/KeA1NoMURqoA/PyTo
X8ZLC/k4Ya0/rzn4Vdf74T2FmuDNuasgfGB42ktVI9YnamMYgAdlHF7TyDG1H9bOPSMETqOHSAvM
qWJtgk4ve8f/H35M3mG/pIbooHLUdL6kWt7DZ6fIeM7DTFMoj9c86TBM4Cky7QXzHrexbVRoOP7Y
btFDUvjNE0CbJyeUAMDxJJkgFrGIuyPtRyTbFo0qEl8L4VljUrKtPtSAVfNo8xt77X3QocajFa7W
qf2zgK9tqAxF+LyTP81zIlBopkMpJb9vAelY8hjhiNJzX8zpqCvUMFq30OdiJMprl8OcpB2AnKIi
EX/IqyfYFkRevasAfLYGsO2eTPaqXqRXJbFsAh6XdGoPdiXr5efWDyfm6FiCQIPxBBRBNqtFnvUd
eb2ovyRQD3M04c5NoyIVFKvkLmLju5VlzkxbgY3u3Vt8ZR1IUz9RC1ad9NuPYPAek/eU434i69X+
X1jTETLNdBuE14+AUezwXMhB/luKdkLESXlbKI4J8QmulHVtrOpqB3eAPDr/9RaeLucFkJzNtgn3
d/sHY0gX+yxUROmn9VDmPfD1ejNKcShOhMlikwvrfOIGQR67JzUXNjtnXC8BTxrfohI6AujqJnh7
byTG+JfAmLMaBY1RCd5MqerwzxwvZoVZjL0vi/G3EkCqrIkjCU2c9TJPJQWaFOtKxfzzd8tWvYkk
gBCl4HHCdbnUlefaY8kCqmfEjI5eFYy6qv3v+I0RDGfPP9jAolrnox/Gn7HhajY+RCFpr/+hdE54
H4M556cEZnAzsGXhGtL1gDxmF2X8pBdTJpWdra2m7nOm+t734BkF8lCE8pZKIZVtP422Dib0KB5L
Qzgk2NIRrItc2k8k1FSIT3ObbndJ4JD9jYFR6s7HV4JQW437DRJIOdt0rR9NmnCZ8smz2qqyf/20
7nDWhAg/MG+SwWmLa+dupI/Xz0pngnKKgWpcfGRlu/Py/RF2uuuYh8XaI9aFxnT3ZrI6duahxWJh
D8GRsuBT+4CcBkRv4/zq+sb0EMEQwaUL1hwtNWPKnfVIko7Hxtb/w0sfL0Uph4kNFI17qwSvf0Uj
p+1uFEQFJEUTzyvKOeU5UXwnCrmfGKpHa0P7jt+ttZvPV9yyRt+bIgSlpXubpQwa4UR90msSSdLN
FLv9jhIZsLkIHJvW8CGeVQHFGaQDV5NTqM98bcLQgRATm6+5dhGStuRj4/H8XG3/tTDMAv2DFf2S
wMZhepwkciUnUW+YYp5hODHi7bSCbgdYaBUd50vI3nUkj3B3CCaq3iALTLzljaLgWEleNbj6xo6/
yh3BJGgA1M1o1KLM/6l4OoHvjWL+DEDPwGIwieSQBJoHkVhVzvwCwfzev1GLgldn/I03yoWV3O7s
D0G7BLbl++xDr2D5LgCcjQ0TmsZbUh6KN11JqF2Y1xR6yUUK+4AfgAzdOQurGFqORwecoIVJI1kW
KMkoIkPmuHTQ+Rf9fwsBm4Tnx7k28bQdxfR11Hr/WkUPNkQxfNMOSkSkt+LlURAdRyWqD0u8GlVa
kN9xUD7811oPd3OiM+jdLCbgoR2ST5LKPa7oxbPfiUW4x/0HBBkg452kd58Jsh3/qQl1jEcxAjIR
EY4IYCiPzdDzCpFOWKQIPFHmuX5ibgtSs86dfXNKZ9EvJpfho/hb/ZsUUfLJWRlK+rxpDdChpucK
S2Y0mmUVi4Yy2Gd/nKRIpVz0QZ8M7142j4StOxnUgCR7PsQ4rP8sEx8Tv1IfkbPBYrRwZxmHgyPa
Uxi5jSQpsiH26EIVyDvUoK1rTBpoa0fELUYdRA3nwUB23zKztUIjFIhgujuoGb6cmdPSc2scHfe9
KWxaPosp4OgfaiKwPanfoHU3bIWiYHr0MUlRMj7l0hvDvVBVTp0ytXe6gTOJq4HMN3E2ZPQjptg9
PeVDcKCAcHRBhw6FC+lqB41JTKGaRvX7GU189dohGoLRqIO3aaXsDYmWdIKu3F9LDBBTmr7lDZRd
RmkMsDyNv49Q0RLsYt1Z6iJyTXHdHWwYRDYjqXlPPLSVzXiyqTeKI2PjfN9meBvAhj3EfN6zHrSQ
C+4iqBuSyjCILCnyg+3Y0aF0IiDkvsuaJ6X6JGs0G0xepZNlDA3FK1YCaX/KyE19kRquSJuLmW9P
GUv7EOfSRKPdyRZYBQJXImZSe8fI7XvmFvPdDV7RsQ2DvOU8KUfaMN4hSxvPlfXXgekRt4Q9PdDO
3suZ/9qu2geAHYQ8BIpqXZRTYFHhzWXmcyZjfMI+CHK7GLgRyjiLjtDjTYaKUWKqXtVoZrDhMQOy
BUAJpijn7LFmtoeGomIl+Wp3FgKuDlJl0ch5XBBCT84NxTrtJd+cZUpO9LpUM/qOxPC6/zY0/nAx
mBTS1Qtlev0X9pP4Jc01EFPWd9r9WShG0HPNQpCPVWzCom9Ru8zdHjExCJb1CRWeQ8e5uLy9RgXX
PDXrJm7p6lbMyZTJO1UrEPMnFZeQShVvhnR0ezbsWZLWlD4cy7ADjeFQDcHpk1jIcjaGh1k4CfVx
UVu/+FGQPmki7JDAy0mfWcp9ZOEyGCC3w+VQYJ50CLMLJDYwJmiOhOTQEmSJcAG75otC8k5JfHB/
s2dsvQz7IwP6rNpz8EcF1uInGBZ1dBSBtNidlVrTe0hrfshw0sQgJF0XFRc9m9sjeLsBV0HhwRSn
u0zH/ZexXdtm+RdJ+3FvQsFgFnb0Rwk6GgJiflw9HxUFkVxxxMGjZ6PIfulVqKf7qhMHgvu3hYxb
Y1iLWmkizlQd+sfBaP2Wjvfpt1L/OE4OG7Ed8MayXnd34SfG/UH06FjbZUoLtWpZCQoY4kmsDRmG
aoCc4g9+O2QhcRP9+6VAa4uQiR3eRngw7fnV6P02KkI8FqX4CrX9vkXAvGNCAgb+tKhA45AydLxm
MtAUtql8MYC6pN68HMQo3pot0CfabAenluV3j8N+9YUOS9uKJz7MWZcNfii29Zu+uyxnDTqlDtCN
IF03NIHHkIp6q3PhtQXXkg2bgjnlczbqyptoR4ckXR5rwiv60cjemXr4k5zCd0C6FZ64SR+Z8FR8
WNVOdytpHX2Fqt6R2xu0eFDtfSWVww1lbRSRtOlWqPh2FYy4SRjLJZcwtctRLZBnBvN9pd5dWHE1
Bx43YUxM7To9oZEnNaL3/M4m1sLpZv26NNz4SpBuufnZ/0P2PZyi2lDGn4+XgatKzjkd+91js2PY
l+YgCIRMDSRItxuRXyCmw6R8exjkuXAnS40HzACodGFtoCFSoMeHPGRXxcgktvNQPO+LMmBd9L1h
43dS4apoiFWjTsQ9Xwwsp1R027psXj2NofGn7I/q8ql0uiUWoFQnPGIyrvk+/bOAWvQ7UT8oPRSw
mpESYY3PMcIAw7w5pplK+o7uT2yr8drvE+JcoKFxa3Je6I0GVF7fGjb5arVYcGxC1j6fuhmiTWAz
Op8ytujI5eUQ3kptGkcKHwDJLkN6GYKObRpNYNOcW1cF+vd2QO3X8o35YPOin+bst6Zk7zNdINxW
nDGy0dxhYrCFRvXg1AnBv0XMVGPo1MPGGnleDxz96zxLK+n2FAJ15HhaV7cJTE6gKqalUjjYTFHa
SaggCbgJhYuFts+q4MvT5i4kyta0H+BZdDSclMFgiEGfBXYYopJH+KhnPRAZJbF9ZX2KN54Oxvip
0WhamYewwVabI4yewMdZvFUgDj7onptDqdAaCb5w7TLwH6UJtGfAiJgTZ/PgXByQu2P551N/PUYr
W8WGMayNebJQoVjJE2bm5fotiEzHXci+E+rpA1G+YyuDz92gTOtuQNIFVmv+KSZN6VY852A9ZTgQ
uE8ACW/TAn3apCyCRBRXAhXhuwUP/idR+khuUGQhQydx74JvqMO1LEx+/IoqEpk8t4xzKtdmb9ND
cz+Gj/EIZX0OHJIvKdFyWIHk8XOXbLGBgvwEJfJwD4brtdrHHvYYCuZrrdzzIodisxecvgXoIvCh
qr1QbunlqGD5a9jHaB+4w4OXDAMQU5zpHF24Lez8PeMX6Vbb5BgEDce3ms9mYVApBe3bbAMH4n54
fo5eg7+iMsu34ZYLkkJUaKC01VSF80GSfqeSIyyRHVrJ5sXW4E+JP9nb71jq/C83ssEOt8aF2zq+
e8+XciqYUQFlPFJWhmhM4KaTnsyJ9leSDEKJmKjUY2KX3IOkX0r8J74BzMDnlEOPL7Xt3DbzHpKb
2poAuGPkCmqFQQ0qlNhUM9hDVQxNawQgsYr+dX3Sp99j39eUyrbxKm0/9cIfxTQrrchOm74WkXM8
qhEZFe4VCj6jm8KXE0c+rnMU/0ITh9jriT3aZGTeB0zNA3zyejGnAUhr0q3Io7Vvob4lIeruDbXU
XgRZ4hNPrhfTbgt5H9Wk+b2RpL+OZ1p2e3YI39lvd+S15aVOB7poCAUGs+1bDH8Z57RXFUB7LJ/z
ikp1qElbogLfmNMnravlLM8wqi/uROXUTjSVjCzDnt4FmTIjAciSvdInxpGt0hypo0vOkpEED3zd
fY3qRpz9JAMZrBe4yRtUuxrYOiWOH05umN5KHXWWJuNjWAI08cfvAxJAWacXkVAAFEv+ca3FfTE0
1AsZSIqEF6mGI+Trteck51yXNL9YAzPHHWEevA93VyQdX0XhQCHLyh1lfYVzQjsTvepkmpp4k/Li
z4Sti52Q00S2RmPtn+l+hjaM9cIaJL06HXFzUEBtKKwQ0ny83BX2MVea/+7tiKIzqCstkntPJVMi
5ooCKsCZv42wiPnjxxBgQU+3Af5owQzZHegFhbth/ezWS7+0+BGbEha35JviqpWODBNPGCSGAYmn
aWJnxl9FC49z/Q+eUHGW4WAYrCuyJ9qvdCE43AdQf5+VJjQq5RunGLz41AsIfj1uNNtP0Xx27EIT
urFh/i99PArGckw2kA8A4gW5O6TexWRkdwhtyiRgPAB+zahykC1FnK7iYEQLc0Pe3bjK994pjPd/
fg67Fqw4ZY8gS8WIl7iAF94dpFwp/zC3jMRJI+0XOw9ORHhqK+xUdV+IwXby6ol/JdNuNHpeIMsq
0oe2e5/nC53b8p07j7TWtr9CfkiEHuf/gzalaLd2VzDiNIpGA/ZW4PlbT7LGEwIVnH7m3P5tLQWr
Z+hg6YsszvG/QKYnUz5kAJ5ouBE39KmdIycrRS72alDFu5cBMi2e6/2qXCl8Afe8NX2mlFFRdpE/
e1CKgeb+QQslH1jAq9sUf5geEHQwFrw8jbI9KlE6iP2LRZtwy8XbLah7rKAcgdsHYixQtsK2FetZ
hwVxH3dT7/3RBfaqeSYdb/cgTsPIHDYV91aydqDonu1Lv46VS0IDJIS3KzyUK0Ohfk8qFY1vVqqr
lYefKOof3hy1aCVLl9e5GwVBmGp8loTzBf+jo27IO7TUdW8dS+m/CBaYLPKKkb9UbpDEYZfK1U1C
Ry0JqjerMQLBYJdzMMAhcn3eSVJn69s1835CLBENxM3FsDEB58olozvyoAdXfttRSyfaQwrJORi2
lHJP/A4xSbpc/KkCnGIAtmMiotuRiIqQea/rzVL/3QMvIv2snUmugqKW4ApcF7+GxewnByP1Wgi2
am1nStm3v4NR4K+qSCqCpThfQPNvuJ2KgIqyCYhC1yU9eQKkyvrHBrFc3RsinT4WK59PH5YmGYpd
GhMKA4rIQfxHCnPPQFKNNzA0lRK5y0o5hUaQ60MgMNmn6/fzHN09covTKnm1dhk+ry21XXCrF9MV
o1382jutrIoUxZaA3zKHlP6WR9R0f8Qw0+oMdWAo4AjEq2n3cJSNvbQSEtYIuxYQ8iIZvnIcoyzU
7Q6K0ZctSOShX2drQEbGAL3SRzlX98RKtv2Vpp6jBZkdwAeE+Kr337xDmnPqxaT7W/rKEi2O8W+v
v1Tfee3WMRMR+/P8/xIcsEuRzvrW/IhqQRhIqzWnRAiMuiyTGi9/wzuygmdtOE5Ct2dXbf7jTG5T
G5y4gDONWCTvx6o/1vToFeZPBlAfPCAjA4UjlVifb37QGwcVay4iVI51sBYp9TLUmy58U9/bXO1b
5XfdGm+QIibsz/5Wp9mEqlULEYVvKIMzW7Q86yDtfnvBKvGb0dpPkp5MhCaYMNnoiBG0FHNcv1Uo
GnC7Cb/U4SKCnZBpHLtYpnD6cq5YXfYoABFhciTyk7nudGrwnnp91zk/LSet3p2rVRxygjDHVep6
MukevJWyCDw75024lqjxPJ2e/atDuOcgk7vpIrD5AfEwzpQ8oCC0Lv/2Keq/HEhsFdjhykZZ5iVp
OpyH+Po+ci+WP8MJ4vhDPocQWPv2E1eNnelwUa83QZDXFGsBqPUpgOsMKux+77uPzZQwH7zYbWqv
tCBgnArcBG8OtKmMwZwtM3vzfosU1geCAwXmQn+Wr3i1zb6FzVteENRD96ao4T1+WOq6ps6jYqWD
/lJgG05u8NBD4KGUIu/ssCbl7DheW0Ek6NivEbK9eyOMYSnuVToX8oTPei6SQbePepQ2MlYCm0eP
gBlwwb/Hoik38T3cogch8QxuRF9WJYYhMMkIqTmLdcH7dcUuQjUQXKKWH5zxq51pQVupX1usGs8B
wh4jzB4wbQLg3wJXpA/O9Gt/0GLNNrfwzYVKyuS8GwAx2amXzkFAhnAAN9OvpsPDRbvSQvk4bHDB
6L+u7fnBcGAXR9hxXEkAJH+69TtZ1Mc5N5uv6OPsV3fGjf3+xm+NE8SXJnhlkz3BXfEgyYCCEx+2
NGY1iJ5uf1VjYDi/pIC81WpO/Ca6YpzbbI42fgkCIOb28jjpfxKAylo+DKISyMqgSI4DkC3kgeTL
4aD4VkzkLzWLgFvchU8DksaVNrhV6va/o1pqq7EbSwwEB8kyCW92qMV3r6ixspUSCH55ZVHtm01c
L300gYBbX0pux5iDsPki43I/8gHCiofl1DpbBuFkF2B4mD3WuPELAruRfmNTCchR107mmbTGQhp1
WrAcDiNK6MeGL0SvMegh7dbHKS4vjtLYibTPJlJTCB8azqzAw3i+ip+VGKW84ix1UQ1PdQFWRzsO
WHV66HCXZOzy0BNnzVHoFPvDBHasNVbCOvDAn3lMfVYpu3dHilHSNeOu79y/uLlhbsX8Bso36KW/
WbhTF83QdHqemlhf0AnGqHPTOMRqqWwKBNo8c0msHocjZru/6/22XTEEIbEEK4cRMcfXxH6AwzVL
BK/zF4S3HAt7ObxXGCldHe0z5exfjfJx2rREwN1h3EB9TcsAAXjBaQraePTIEOwI5vNram5HbcIV
6HjYPDP2oelHlu8Jl9emKcexGfP9FhXdHnyPNavDq30uQTl1ssXuE2uwXRss4TzfsvjY2nOae6BP
fkqWC+c4LYeLvIc0yyL5Id7gmTzmNWg+j8WcQQDla4Kuu+Bpbd8sB9xByspkWPvb7wW+dRrtLIJc
fcqO9wWBOAPp
`pragma protect end_protected
