module gw_gao(
    ready_c,
    \data_out0[15] ,
    \data_out0[14] ,
    \data_out0[13] ,
    \data_out0[12] ,
    \data_out0[11] ,
    \data_out0[10] ,
    \data_out0[9] ,
    \data_out0[8] ,
    \data_out0[7] ,
    \data_out0[6] ,
    \data_out0[5] ,
    \data_out0[4] ,
    \data_out0[3] ,
    \data_out0[2] ,
    \data_out0[1] ,
    \data_out0[0] ,
    \data_out1[15] ,
    \data_out1[14] ,
    \data_out1[13] ,
    \data_out1[12] ,
    \data_out1[11] ,
    \data_out1[10] ,
    \data_out1[9] ,
    \data_out1[8] ,
    \data_out1[7] ,
    \data_out1[6] ,
    \data_out1[5] ,
    \data_out1[4] ,
    \data_out1[3] ,
    \data_out1[2] ,
    \data_out1[1] ,
    \data_out1[0] ,
    \data_out2[15] ,
    \data_out2[14] ,
    \data_out2[13] ,
    \data_out2[12] ,
    \data_out2[11] ,
    \data_out2[10] ,
    \data_out2[9] ,
    \data_out2[8] ,
    \data_out2[7] ,
    \data_out2[6] ,
    \data_out2[5] ,
    \data_out2[4] ,
    \data_out2[3] ,
    \data_out2[2] ,
    \data_out2[1] ,
    \data_out2[0] ,
    \data_out3[15] ,
    \data_out3[14] ,
    \data_out3[13] ,
    \data_out3[12] ,
    \data_out3[11] ,
    \data_out3[10] ,
    \data_out3[9] ,
    \data_out3[8] ,
    \data_out3[7] ,
    \data_out3[6] ,
    \data_out3[5] ,
    \data_out3[4] ,
    \data_out3[3] ,
    \data_out3[2] ,
    \data_out3[1] ,
    \data_out3[0] ,
    clk_byte_out,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input ready_c;
input \data_out0[15] ;
input \data_out0[14] ;
input \data_out0[13] ;
input \data_out0[12] ;
input \data_out0[11] ;
input \data_out0[10] ;
input \data_out0[9] ;
input \data_out0[8] ;
input \data_out0[7] ;
input \data_out0[6] ;
input \data_out0[5] ;
input \data_out0[4] ;
input \data_out0[3] ;
input \data_out0[2] ;
input \data_out0[1] ;
input \data_out0[0] ;
input \data_out1[15] ;
input \data_out1[14] ;
input \data_out1[13] ;
input \data_out1[12] ;
input \data_out1[11] ;
input \data_out1[10] ;
input \data_out1[9] ;
input \data_out1[8] ;
input \data_out1[7] ;
input \data_out1[6] ;
input \data_out1[5] ;
input \data_out1[4] ;
input \data_out1[3] ;
input \data_out1[2] ;
input \data_out1[1] ;
input \data_out1[0] ;
input \data_out2[15] ;
input \data_out2[14] ;
input \data_out2[13] ;
input \data_out2[12] ;
input \data_out2[11] ;
input \data_out2[10] ;
input \data_out2[9] ;
input \data_out2[8] ;
input \data_out2[7] ;
input \data_out2[6] ;
input \data_out2[5] ;
input \data_out2[4] ;
input \data_out2[3] ;
input \data_out2[2] ;
input \data_out2[1] ;
input \data_out2[0] ;
input \data_out3[15] ;
input \data_out3[14] ;
input \data_out3[13] ;
input \data_out3[12] ;
input \data_out3[11] ;
input \data_out3[10] ;
input \data_out3[9] ;
input \data_out3[8] ;
input \data_out3[7] ;
input \data_out3[6] ;
input \data_out3[5] ;
input \data_out3[4] ;
input \data_out3[3] ;
input \data_out3[2] ;
input \data_out3[1] ;
input \data_out3[0] ;
input clk_byte_out;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire ready_c;
wire \data_out0[15] ;
wire \data_out0[14] ;
wire \data_out0[13] ;
wire \data_out0[12] ;
wire \data_out0[11] ;
wire \data_out0[10] ;
wire \data_out0[9] ;
wire \data_out0[8] ;
wire \data_out0[7] ;
wire \data_out0[6] ;
wire \data_out0[5] ;
wire \data_out0[4] ;
wire \data_out0[3] ;
wire \data_out0[2] ;
wire \data_out0[1] ;
wire \data_out0[0] ;
wire \data_out1[15] ;
wire \data_out1[14] ;
wire \data_out1[13] ;
wire \data_out1[12] ;
wire \data_out1[11] ;
wire \data_out1[10] ;
wire \data_out1[9] ;
wire \data_out1[8] ;
wire \data_out1[7] ;
wire \data_out1[6] ;
wire \data_out1[5] ;
wire \data_out1[4] ;
wire \data_out1[3] ;
wire \data_out1[2] ;
wire \data_out1[1] ;
wire \data_out1[0] ;
wire \data_out2[15] ;
wire \data_out2[14] ;
wire \data_out2[13] ;
wire \data_out2[12] ;
wire \data_out2[11] ;
wire \data_out2[10] ;
wire \data_out2[9] ;
wire \data_out2[8] ;
wire \data_out2[7] ;
wire \data_out2[6] ;
wire \data_out2[5] ;
wire \data_out2[4] ;
wire \data_out2[3] ;
wire \data_out2[2] ;
wire \data_out2[1] ;
wire \data_out2[0] ;
wire \data_out3[15] ;
wire \data_out3[14] ;
wire \data_out3[13] ;
wire \data_out3[12] ;
wire \data_out3[11] ;
wire \data_out3[10] ;
wire \data_out3[9] ;
wire \data_out3[8] ;
wire \data_out3[7] ;
wire \data_out3[6] ;
wire \data_out3[5] ;
wire \data_out3[4] ;
wire \data_out3[3] ;
wire \data_out3[2] ;
wire \data_out3[1] ;
wire \data_out3[0] ;
wire clk_byte_out;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;
wire tdo_er2;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(tdo_er2)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i(ready_c),
    .data_i({ready_c,\data_out0[15] ,\data_out0[14] ,\data_out0[13] ,\data_out0[12] ,\data_out0[11] ,\data_out0[10] ,\data_out0[9] ,\data_out0[8] ,\data_out0[7] ,\data_out0[6] ,\data_out0[5] ,\data_out0[4] ,\data_out0[3] ,\data_out0[2] ,\data_out0[1] ,\data_out0[0] ,\data_out1[15] ,\data_out1[14] ,\data_out1[13] ,\data_out1[12] ,\data_out1[11] ,\data_out1[10] ,\data_out1[9] ,\data_out1[8] ,\data_out1[7] ,\data_out1[6] ,\data_out1[5] ,\data_out1[4] ,\data_out1[3] ,\data_out1[2] ,\data_out1[1] ,\data_out1[0] ,\data_out2[15] ,\data_out2[14] ,\data_out2[13] ,\data_out2[12] ,\data_out2[11] ,\data_out2[10] ,\data_out2[9] ,\data_out2[8] ,\data_out2[7] ,\data_out2[6] ,\data_out2[5] ,\data_out2[4] ,\data_out2[3] ,\data_out2[2] ,\data_out2[1] ,\data_out2[0] ,\data_out3[15] ,\data_out3[14] ,\data_out3[13] ,\data_out3[12] ,\data_out3[11] ,\data_out3[10] ,\data_out3[9] ,\data_out3[8] ,\data_out3[7] ,\data_out3[6] ,\data_out3[5] ,\data_out3[4] ,\data_out3[3] ,\data_out3[2] ,\data_out3[1] ,\data_out3[0] }),
    .clk_i(clk_byte_out)
);

endmodule
//
// Written by Synplify Pro 
// Product Version "P-2019.03G-1-Beta1"
// Program "Synplify Pro", Mapper "mapgw2019q1p1, Build 007R"
// Thu Mar 26 10:12:30 2020
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\e:\gowin\gowin_v1.9.3beta_37257_win\synplifypro\lib\generic\gw1n.v "
// file 1 "\e:\gowin\gowin_v1.9.3beta_37257_win\synplifypro\lib\vlog\hypermods.v "
// file 2 "\e:\gowin\gowin_v1.9.3beta_37257_win\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\e:\gowin\gowin_v1.9.3beta_37257_win\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\e:\gowin\gowin_v1.9.3beta_37257_win\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\e:\gowin_work\ip_design\mipi\mipi_release_case\mipi_dphy_reference_design\mipi_refdesign\temp\gao\ao_control\gw_con_parameter.v "
// file 6 "\e:\gowin_work\ip_design\mipi\mipi_release_case\mipi_dphy_reference_design\mipi_refdesign\temp\gao\ao_control\gw_con_top_define.v "
// file 7 "\e:\gowin\gowin_v1.9.3beta_37257_win\ide\data\ipcores\gao\gw_con\gw_con_top.v "
// file 8 "\e:\gowin\gowin_v1.9.3beta_37257_win\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
nGQjNTRggZWOT6sWc6oyraDUFLfWAO/HbLF6wXbCqXPNp9WCDJpv1rHVczOIVgncR/b0+UeSwebZ
OxlPzCeuO1qPl8FPTKiUyycPd+J0aSTr5vl+//g43DlAnrAZWpp+9NwkyX7Tl4KQV38q+/ZFnqAd
fKrxDpwkhDu4v9GmdKTtVryneeZJtk+qfqQLeux8ui4DI7WokBCiLCcnunBZc7zPDJ4RNHhhj/d6
kphLiA+2e7BZhQi3+S17OFvZZeAZqB9QHyWn8tsgCw/p96pTPtatJ/h1TGMYgxgbBmCeWweLMmye
bCwg5pbhghYptD2zVIQFJWuiylXMfypQ3ZpFdA==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
x5gHfLwQ9h6IkqXYFQsKYOoMTbgAOviKZwc0Vf339pYT772gCzJCT3UDF+YsUsYbK+Pq7BKRT6Uf
HBulNYuf7y+Ku9k8h5gb4vT0dUa4DG8OSdHb7R0AC/h0AeBTlns2hBJ4OSQGxyyNBp2s9HonSdOM
8ZWZFAphVVtPxikUpfU8q9qzyHTb9jMLF3VfqHt1hy3qcsmu5t+UPmv9c2zjTl4NXRMUl5483dXo
fMq4baFS/ju/wiHFuRhteazMg0mM6BfGhtM2aDlFaVzlnFbwItgar6Mu4Fk1u80ynR+wqXfj4ur2
96zU62Pm3UBbG8dYUGOAgfAhYDkhAs6USGbytQ==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7104)
`pragma protect data_block
S64wz9lq30aLaC+kL/X10osfDUSymmrQf6hdQCYuLnmlW6w0Fzin4aO0g/WUobnGsoCOY7+vwaK7
shINCGen4o92p7HrSWBdN+5Baowett5dwKHQqJmKXDf8kRu2EUM6L5usvI7gmjwb0Oqr0AOxGdMA
IEt240OIHMHC5+4DWcK1R5uW4oisAZTZ0NJomTQDaMYTf0vbCXRvBfHpZ4l5DtYYykQ+1wrCdaX8
sSH+7Kja8QmLHvKxnpa8f5JIgVG/ucAiaLjJCwWMxb9Jgg651lo4it+/5Tpuo5y2qsnz4H1JMNUn
Uj2Wb4mlOEYAAuxfOQgISpA8CPBcEc7sbHGRaiqACMoKpmzuzNxNUD8P5cv6ovUqQfJUioqy8RZU
ncsdMPHyh5mNATv+rgnC5o/KV93EFFByE293XvqXEYEjt9+B0tjML3MngPfTex/cJ2bRYI1Y29hm
XTL62PjJKbMzmK9NpFeIkHzsZDbc2u2z/BIavl6tVtDLm+SAcnppavWyK/5wQreqZ2yB53u9z2o8
LprLjQ9sr4VB4syjJwQmDoIF3R2IbM/QcfbvefBq4dq5wIAzfUOIsG7ArZLpKq5bpD2Zb8A9OHiX
uvKXXGCAt2zRRcVLod4NupUa6X2EHnU26zdjJmoMtd40HPn4cS1oNYsj8oDgnMRuf/Usf2EPCPzZ
zBwI1jWvbx/LDqAKeiJy5p6Z3ppYHfexLl4KVFJwvZN/UAIWIEdE4gMnasijR0V/X7zNIff2Z+mg
Vst3itLdrWLhIpU72gmh+FTfXmgP5G0QzeUXu+8N1eSeRol7/A0ii/TmT6olTEgp5qz99PEILD9D
dwbTqx6rbR/vbvZYn5A6MKVaJHf1Cf2AGsVHwSde1kyO3hEKtQ4r9nRWUIdDLZuN0jDbKAOGjSOj
cKQrNjYtn3fCdAE+vAydqBHJo0aNdCmOVR4Q2pRU6nYrm/btQlG2q7hLFtC/KPp2DUkDmxN8r+5B
jtXBUi4kv0tFiBkb0PSxuTRWBbmxgMHvu2TByRH6BUq6yGS45JSdbjpP0iYwguTga9uQlQJseJvN
j15bPLNnu23qzXFj4YABLhVMn3u2NXCFJtuYMqFQMW1J4orX1gR/oDz9x64hSD6+sdyOMqp9gEDe
0WZRRJAd6GzrJiG2fvPM1m81XHvAT/TIg9osTlKtlSzXzVuRYotP/nj+sMrIXuurrsc1pfn7ea2B
ISrslDG0drHlU2Z8sJzhGbASHunb/c6FDO3xa0eSWtFJY0Zhrrea3oMJs//S0utiBr2gbKpvy9fe
8P5r7IOy8zteMADi5GQL4tpxJV7mLmxV5wMl6chKfGEa3EQLt2ewF8lwfO4MxsGevQfwzpyEMxeP
lSwplNFiJcp0Xv6tqh8XEID1y/HeVvvgJ9GqNvQp7IRjtyofC5cnYhdVZgSfZnsxVLMI9XrEy4F7
1kcZlF9qPaqvan0/v2PAvQNTE4Aky7dcvYIlwEPyugt1oVg58aKh2BmQeOJC2BMlk3I2WanCtp91
ZnKNuFzPrfhXXPj2wxHeiSrocPg+CXUwYn6Lh9ZP1CSTIgcTSTO7Je36R0cteVIP6MC0dl3CNe3+
ehIH5ri8Mzq5h7hYZ5xPN5SxlC6R8ztqEmHBI2n4ocW6PoUJ08k73moWX1fffyHI/8+PJXUZQXcy
i/QOTYTMWNe501G7rJyE+LyScYgUc/omd52qfR8yReR2emmNkCCfpMAwNRuD+Obrm6vgnVLD50LC
aja4BCvetXXvPTbxgWKx1O7Rb0rcq//qtTkZP9zmzoslA8sCxkHWScRmmu6PSlJil29H3gdvNnRE
2NPXv72u0lDva5U33a2Jnru37uCEX/uUz0xz/bzqIOf6UaR2Km1sgblMqE3ShRNeQjQIuWnOH1Zn
f9Cq+UJBPgdeVfVLbIWLKT5i336m7o9HlwZplVN7eWrhxkYYoz/R/oozCpwRu0QvpA5o3zE7v52s
WIBoKbw4KO3Z8tCfCgBZ1y2bYb32vB7HINbQx2k5MJ6kxmNJKYPrxeqku7ISrxm9ovUD7ZsXWpZd
oewJ44kZko+tVZFoLxkhKeUKsOVKR4+Ew2XtMNbgOlRdz+jrMobvgMRKr0/AmXYkZCtt953ftRFz
D0IRZcmDDH89fVuKKj107QAqMuHwQrByKg0/PGinO0F9HhIhrhys76y1RNOmtZ1aa1W8/wX1Q6f8
vN7j6FzQOm4zSeGTjB0eFw4I8VtnVnU6X64M+KcatrhMhjU5ksH7weN596vjXsApbnjFkZ+bQIuh
+7lAQkAJTrAiA9vzFZPJ9mrIxf1k4By/+RRZplp4ECFu5Yzf5D0iwm4jqHmbUdke8LPcjZ8rmgav
/hD6yMURUV/NGEJN3DGT9CO9W0MY4ZFVbIQ8oUFlw9qaytzJF3D6GUEFf8n8s7ZLMkjcLCyouKYS
HsYIdM+JJfEhsw/IFdI+vy8rjjuY6JzqFy5/C7kwTjnMCWWFsx+IQy6kIYNJKKqdyH4A0fL+IWgj
Wk5ccaiB8Fc5kP140Yf92n5SPBGntrZ+z0OR9BA44ousRetZ2iPoJubaJpLqJqITXanOwv+GaYE2
xApaKCCpBpXaWka3ltAXvIX+J8y1uDraEF6X/qElfK/QUAlCItZzzxDjuWjKK8V8hcjsHCRIl7YS
wCFkKNjk5B+NtxB7gYGmfUEDxrN3rlhj+9591269ETb6mGGlUG3fk1PLQu4qbXt011X1+Tui3j4j
t+iahFSKekuQP1mvV2eRD4wxiIaUK7ZOTHLdCOSGulU3N+EdCyMizUnXj0ROIu+4/g/topa2fAly
82E39Ai8flzWfclKLaiPeSI6f4JOuMjPs9rZ7bikdDZqVOm3Uq0AX0dQwQoWl/H7e9jWg/fXRLNg
1ha6u/xqwBb2vcrJMgxzW+bfomcC/qDenBNxlMXMtuJAw8xgBt4/6pOD+N02tMcvfNyjrQBlCpEJ
r2XfbqlT7ZB96dE5qtvq7eEbkNCyjNO/psoxV6y9U90VEz0oXTG2cq+eNZSikQICFP8ge4rDenfW
asHDeBLqMvP+bFVDtTZ4sK5dQC7DpHAvdAzD3+nSNyViYnY7ZR4nqcyeBMsW8yV+xQ5xyaZqFNNZ
84llEyWvNtn2+0j8ox5wU+g1Ozg+bivHS/Ov43A9Q8en+4TX9Q7et225rLDi2N8yt2yWrBVrJOkC
sIsxjiPMXSyFziIytWlSTNFOZBecpQJuVdQMxitP+8KDPMr8cwXlAGimCffnTjbS/2AxVF578yj2
zAIiwgVzrTwoKdO5qp5bk/7Qxm0RHiu08lHOHmH6a2epkeywUUp83PnHICHwIh/6l5FWN4D4avbe
8eh1DaA9xSr2w7MEMxGcc+GaU7rYw2YuHDhnPtViskDE+g61yQNpRER6R3C7H3czbroSXZ01PvvO
uTbnB51sRBzatXs2XAfKB2BOtOK0xfKrZb7TuyiKjjZjZRIlbjWE+3OKZwHYrYuIwLXjNfzFww0A
IaM8zPtaPERVSLkWzuli/hREbu9QV3/xinws1KQYARjR4mimZy8hmM/nqWb4OF7Cs/FBMU3CDJ+y
IfRTlBwn6fKr6C3IjBUd5nUDVhCXd9ZD1BDFztCwEWRntDyTI4et1SEkmcgGuMPYIWpR10r4+hkT
oWyg70oE3jADAbMBxP/rEq03S8do2pnaR8L2YK2AaCyEgo+jDZtKD0TxTBhWHJinpeQDLdKMrJFP
FrkZkzXMqfucEeVbtlvDI3H7GLNgJrPmuhq8zKjcCmDW+gPHFrSxtqAvUmkurh/vEiR/SDH771ri
qtIcbxIbuSF77nUUKPLNnW7aBU3c4NSkq6rWH9BixiIPoQII9GizoYmUKJ/X5p7yWotFME1eEQ9j
o1wtUyT09BdG34lvecbVMfIlmYCq3OjDNPuFgte6rnQtlaNBVEIqP2zQQQiA+j2P5e9oN/fIy97n
QFbcPFkh4duzUZNsLrzqlED4xklpzuWfCMTRSzlYWSPYW+HZ8sQ5r0Vtppdw0NRJYGy0S9o2dMRg
MvR3r0AUi6ujiORnjUk1DAqJBF5bFT68UWKMAjhHOx+4Lppz+4/KXQelsdEIKh7R0eI3edF/CXLO
/cxV4ClX4cGi+jKbAjxPkO4phmx2D0jtgQAE7Lvq8xwGVI8D9uuNccq+EqxEYyqkYCxb3PCzcUAG
aCkBvx4CLL6GMxg49LSCdY+8ZBoiNLriEyQ94IDYMTXaHH80Se7FF5ixNjcgfthf9t21lzxPG7gT
QKipnExuDEOc6Gnu6ePN8g2LI8GM2WZ0bHZ/Fo7KJqlUtSDzM/ikrBfjR95uWeVcWQoQ14lN5pY3
80eBTGp8wOpksbiYZVYieL8nfoUzIJcLN33T09lfaxL+ugRLh5JG8POgZ9UvXO09yjUgvV6evL9d
4xxf1yAngW+Cx2oEuIfJks62f2UM7HGk5BH5YWTM29p7rCZLUinUNoRSrBe/drElyHxZ7AcYqghQ
iQ25iPkCc2jkP106ntmjrvDekZjWCiOuq10UHPG3nwIVILyPsSPRXzYBx66DUkqmHr1ftiTWzQ0Q
/dEhxdrOFPd8G0OkI6Ywdy/hodRpGgv0GWsdESUMzKvWHocINNOYJdn+JIEhdNKjhytuhkdn6ITv
l3syCJWMnZMQwG0QkgvVIymbJZGXlOUtBPGnVNoXjH9S0nXKcp8x5aweNtIHWwZAbjk1j90KUITC
TS1F6ojQfJPtQVO5n1oH5Pebnw+oJK/Ut3mJTj9H3NXlFkdeYFlI4PIiJkbRZSDgidznB/2xyEhC
KO31MVeIkWCxG63UMU+me5ljBDt802bdj5Rwp3yZC25JdddSOrw1mZ7Zx4+H6NA5Rrh9gaIqm3OI
wiJRnCC3kcl0BpdTRhAhp5Upex7zY45MWd+AWqE0WZgw07eF4q3+kNvwplt/JNf9gJu/R0GiP/7c
2AxHwKkiFXoYlcekSgYgITKi9gicgO9mzVerDu9IFK5MrMwwJElKmLLXVqQMZh6NRbzMxZb8CJy+
kblhwgtyOZ/0FlgXDYn3ZDYcyU008cXwB9UvCagjfLMYCJta+Uaoi9/9E2Ch7QYKa8sipLfZdNv6
K6MlqPp0bBl72MRwpOjkRdghaxWR7+DKDnjtW5v1XWXGI+5OgH2LYwoWIYHIt+VrycfdGKpbMhTT
BrRk1aeKvFUE5IPn0IZQL6xhKKEmaoz0j1lclKh/j0he/gz1wZ12n9Ke3tyebTHMpDrN5kujVJDl
te1O05n6pu4w7uwPhiU5Im9VVZ5do6I2e1Vk7J3VOrUMfKftmQ3NToLCK3TjcS2ePO7J9F6T5Z9m
tz2M/XX/T8HfGTmjE61f25+3VeYR/OP2JgxVcH5595dyO3AHK7q3tSdZgPwcsk/hOQq8pTivpTkM
4Ye/Iqzd0Rb3XWHa6snNjCOqiTqYYXP2UxYzvrDnf2KS2a9Bg46nEFdA0m8eiXmcbiTGAgqn1JKk
KRhmqOs7G2pGj3wCZBl0R7QChT37/N/oN5YVawhlJbIluaNH/kIv+Q13wbO9Ea/4HP6lURoFUg52
qO3XS79/wOQesMjUgxQVxMMUI1eIlRnhZGs/vuLJF2kmIS9QK1Klvu7jjmOUHlxB7grS9CHB2KAL
Sc9BwZjxp+v316sq8+98qI5nXKErU2vTUod9/IiZ7yNmY5DGqxqkuqfhtX2FzWfksUsl+B30mRrE
+QxYKaclQUGNXoqjm3xMVVBPOt6ZbcTU+pjPcgkIkyAhMlXE9AI7CkdNG+Tsy7FQzUAIWapQPkQY
n0jyM3+PlV0BMBJGdkIDPvO+ybEbmKhbdnQeRTLaQa5hGdnZ6EMU3y6BQaYIc9jhxfZAruYGDijv
5syCVCLQHAzuRWFcid02IX9ihcxvoe5MYiv3IOw5RnTxUT7uR41vmE8xDytgZtyAw9BwX8492dcC
gSo0RgyonfSEf9W9KGAZlnCTSGdl1viwNCFnWcCY0EB+1MOhSrtfMJiFGPCdnNfa9jPwkStwqW8A
iBkB9E/B4zHCgwrnF0GVMvXqZXnbInVHUJUeB7H66d2y7uwLDtmTKheVWBZELgHF4QxxOuOqjw9v
0BHLZAPYJjwNAWhk4DnxXKRWrDmIbvVZi5J9cahi0Z76snKq5VuJXmg3Hvn3iquNkPOslSLmIlYu
7EQLD4yz5nC5knqZBKX2Iasp1JOE+KGHIhRmlhgRz1j0UGI2FxcxXAZBFe7lBCB6DLlALHRjDMA7
kwunzjIfrenajN4X8OjxpIHxgkKyUrhzsDQDCVSwvihs/cxwPPXrcjpwO8pwpWLIoyQ07D74zW7W
4Xtvz9mQDNGNv5t0S6hnNtHD0p89XBYg/jW/dPTemfD4FqVFU7W1lAhKhR7x0iS+I+Mv0RkY70Q8
V+eSpfYz+vApl9vHY/1kDqW6lO6sCawllgMTR4YPY32/kzQfPku429SQFZepGe/VgaWpu7WMlB/7
ggjYuspkN0CXproD6TTH4Aqgow8txDk02Vg2wI+joePmS+oeVhFTxNG+Nrs0It5I5O3Jj5h3Aznk
bSjboXMbf1wdwL7Tt60X0Ami6t0QVrYKCxEVM86Xo8tK1K1JDGwT56vV7mPC2TBuk/FYhFlttdC7
EmwIvsqvSa0ZCuMsGU7OsvdwnEBPl6JC+12fQUojHVNr3NX2ge7fWRySynWwehZviYk3E+8dRnSY
uVxcGJj1gpmBBlVaXI1rrNFpSQyZovEMo6YHtsnSNDBdw1wC5hOSLTDVgO9FFBgDn8qAzZhAUF4s
TlZJ/kDg03ff3kju9td8fqHStgXhe8606NfwYPagCrievfbeN0Omd0IpuoeyfyvjzJRLbfU+0TRp
dffgRTBU2q6CxGeJB9YKJarfPTu8MVd5YQrxBuwU21VLCBdJsTyOskaCgyRKyRtL7gvFDdpPhXBA
vQoyXlsRBi82LFlsh3lYn3uQ3Knfj8paTxKb8IpLeEsB8BrK2qyPd6koRSnNNkZla5dNCnnx+u4B
GfSj27uD0+hbcCl+0gib0q232ueWUI2csgyNNKlmKkI0YYy3zMLSvhYSsuX/9uJFd37HoA6lMwho
SXel3kNXNBT/NKq8UHsh+WCfS/DG7dtgR1gT8qx5fG7jvnkyh9tvI5RrqhVcCiwrHOpNe73zXzH6
yzDtESL/55w3BhjuXcdlB4s/+v46azuJEPFdFuQzQfgg65zQI+NncX7KPynxJ1UWVzCrlOib8XjK
7C11ON1/NWBSpORI8hnITmzSZ1zzeVZxjXBn90jtMZZPpk5gtgsHX8BHRIOUSGa7IfX0K4BGdSW+
2Hhzk4wz6+CUr2bgVLqPfbjmvaauSzZjMHaG5qoVWVnsXo6/qiOrZ7eENmsTlki8wanOs6dgYfj0
vp1H4FGqj+mDcNI63JXSMZaa88DsNabqS2w5ipuYGgGxwfreVwjzJzJRPYqxeehXAkdF5ZBRTcvV
QWkXHgsqRSXyRoznuokAvcHJ+JZf35Cw1S4AvL9bTLk5YT/c6sz4A+H11Gj2YVZ7hJ5Wb3/nn+b9
Sc2VYSORZV6KkZkhysOrUo9xF4NmJqvNMfdiizik+YTUQUYLJC604jflRFcJ0KHEQyevJQbpm9Kt
jmqPArFRgU4oUCejVugs7ej0lJA582IBQWT+TGp9/DY1G1odWVXL+UK7dm3Hup9cQwAgv4/sd4bw
9H4hWowE/BFhR/8i8EnK2+gkGNmEvmqxs6mAJDoj1odVZ2sTtoTAt+M68FTruJpQsUxXeNdSkaeF
TPvrNsjqI63/OAjWnVPvFMts4Ay+DfFyLzf2xOoUZgdBo9tQqleA/Azac+VvEVr3+PdW9MNiaH7h
PQiWyzHUUC3fnsejIk5/xXo/pttJrxh1HI7iS0IdMmkkY8MevfzapSMHIeZFZwaZxlvUVeb0rLbh
scepHjwS/TS+q+/KAgsgPYgI+Ok/feY6hPEnRRI5Wj4dfshbDrK7yFgVIJOgwC9xTmfiqh8gnbaH
TFvy3PdHKIZ4tBR/tGVFV7FKFhVNaSHvtedKfHUMnqZ5WzEGAHdrnNwm3UmK6OzG8R2HE7P3P00F
pPnJppATbWaddStqZWc0l+uigR1XvKoUmPRIO34kwcka17ByPa7TLeb5LY/pYJcTO5ImfVnnRZQF
UDFU9Tusr0m16oDdJLLfRLAFzyx+Hv3EdRfOgbC87mW59a1XQ25jKWCvxEZrd8DTeltX0AFWrxFP
X0l/gfSoHnaGDREhbpBtlUC1DF7yn1vLII9QnUTCSR9xkt95Og/nQjO56Q/cUU2TDDgEmHmOjlJp
9aj3RNmlScim4Gg14ob4xofrLVMBJ/H7HJhzCm9Ptp6jsVu7/dDcgk0zMDMpj9mpVwXo4on5WY78
TcHH23RdU2Ucx4U2RRUB7mJHa6y41xQlt88HUVtW2ysFmRocgOBK8ealkE/DRiIuogBfpZzxZ5Wd
SbwxrghO0HEU5qfQUekWIUbRt7NHpMk0GwtYYkONwvHMUI66ZxMlxBPi+Uj6vnHnACjYI7c9pb4g
2UyR7abHkXDe7SmAuygabZHa894hnw/10HzwRIGA0lV0vDjHjZgf/zuMdADV4Ts0ifnkdfx2sm5Y
3tPumtL9qd+1IsoYbB0bogFkxdxhoMt+gDvewCusRk1fmVcKmAm7LgIzaFnJo3TQB2Ik2iU7BggC
0d5CuKCXPFsxLz77iQ0dbHD/KHB/zGyk1xF3Wdq+Whnok2M0wK9M5nyNr+/eEHPIxG4PykGBOS+T
ezvSwkFw5RPhhhdHWVM9ntOBvcKn9KJxZ3Hw8+ntV1i4ul3Z5U8nFc6TGPaPWZhoQGBsQ+GjJfZO
FXe3pje6w7UOr2CL9NSpa194Ew9wxMnavCrl/2e78AKhITDkJnxklMWaRBFmNb6FHWmYm8eicm9T
/iF8rzYkqF2rna+nf/SZAlPocDJZGrJvZR73D2veuxzEfKqw0vAmXSpgCZvIMVqd1i0+djOc1+1m
bdcsXMG8Hh9hjpNGlnEDgQvpDQlUSBcvD1E1tTv5re1x43pIqQ8cLdTrNWh60b2rdlgfYJDk2nHk
VTeY5uQoMAIEqiLbdpwniBkZeXEsHcg4ogmygwk7SDUxVttHiI0wCfgpE+5CY5kOq6rq+nN+963x
fnZSUlt58fHSfkbEDXtjzqfj1xMdt9vFcjZ7JraFozqSYzjzcJEMSR7DsulKIMTofMx6TYVSTpl1
VdrBT/GM9FtMUfjMKjJKtzKaKx+ogriIE6/7zzS06nSKPqWcwzD1qgqAUDSiupXxHn09RiIybw11
T6LUDnrSK5GbcIHnMlsSjEHgYhgc1/YziRRSrDXabhDgkfsHWF+Ti38hov8C1z8nABB3ULae0pRb
U77cmqAZ0y0zSfp6UAQmQ9DP2L69WerQVaVbLAAo8QK9DFC+9ZPP0C/MvJC8iv6CXEglAdsQLTzW
zAmm1Ahe07fWA5eChI/RwnikMciJqwEL/GY0tJ6sGoeCJQu3
`pragma protect end_protected
//
// Written by Synplify Pro 
// Product Version "P-2019.03G-1-Beta1"
// Program "Synplify Pro", Mapper "mapgw2019q1p1, Build 007R"
// Thu Mar 26 10:13:24 2020
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\e:\gowin\gowin_v1.9.3beta_37257_win\synplifypro\lib\generic\gw1n.v "
// file 1 "\e:\gowin\gowin_v1.9.3beta_37257_win\synplifypro\lib\vlog\hypermods.v "
// file 2 "\e:\gowin\gowin_v1.9.3beta_37257_win\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\e:\gowin\gowin_v1.9.3beta_37257_win\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\e:\gowin\gowin_v1.9.3beta_37257_win\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\e:\gowin_work\ip_design\mipi\mipi_release_case\mipi_dphy_reference_design\mipi_refdesign\temp\gao\ao_0\gw_ao_parameter.v "
// file 6 "\e:\gowin_work\ip_design\mipi\mipi_release_case\mipi_dphy_reference_design\mipi_refdesign\temp\gao\ao_0\gw_ao_top_define.v "
// file 7 "\e:\gowin_work\ip_design\mipi\mipi_release_case\mipi_dphy_reference_design\mipi_refdesign\temp\gao\ao_0\gw_ao_expression.v "
// file 8 "\e:\gowin\gowin_v1.9.3beta_37257_win\ide\data\ipcores\gao\gw_ao_0\gw_ao_crc32.v "
// file 9 "\e:\gowin\gowin_v1.9.3beta_37257_win\ide\data\ipcores\gao\gw_ao_0\gw_ao_define.v "
// file 10 "\e:\gowin\gowin_v1.9.3beta_37257_win\ide\data\ipcores\gao\gw_ao_0\gw_ao_match.v "
// file 11 "\e:\gowin\gowin_v1.9.3beta_37257_win\ide\data\ipcores\gao\gw_ao_0\gw_ao_mem_ctrl.v "
// file 12 "\e:\gowin\gowin_v1.9.3beta_37257_win\ide\data\ipcores\gao\gw_ao_0\gw_ao_top.v "
// file 13 "\e:\gowin\gowin_v1.9.3beta_37257_win\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
DI4rXVSqQQakdxUiFbNMpUcFqLtxiH/v9VC2fotO6RT5oJx4ujfd+d8ntglwi9SznfUhuCDdANfH
XYMgV7tqilOQ2ZawjyjFzCrZ5SPXrGgsruT0nRljnPbi6qkiFtugOcQTRLawx9T7//cBM+KloXTA
NW5UEesUVY6XIevfIUZGJ1ure5Ny3juAG8DwrfgVKoVsVbpFHGqkn14/CuCrPfgd3cNIeMnz2tdU
fIIQcJuw7/y7oxsPIHnSNjduB2VlABUbTul3/U+MLlIz6QrQXnGGd0gsk0VzmjNw5t92AUKNXFJQ
KgZfLCLpjgQ/ZbGsMSNTxIFdLQdlxHMJmC0vaQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
BJq830S/kOcQBA2JJ2q4S6I8jB9jjQ+2w4M1vD4Tqw23sKPDOhifxjr0/o3W8kskkjrPH5ExmJnx
4+Ax8NsC3/y94RfnMYtaR48dVDd/uZPC+H97z8xQbMlRtAPIPBxmvbm2XF9esKwvNQk33qXslMT6
Af5S+VRtkbzP466p8XNJQwyztsU9oaM7FXV1jV3HosbJuRzcKVPEOmo4Dn/DOSxaP8rd5LPjoLqS
+itgiiOB0/sBM3oF4lMqNh90Lt7h7dN75Xc5z0AOiCtIi7ReGbnoPIxpLrTX3YY2f7/TaNJjwe2m
A2muDv33kmPJYj0Qn1mVE7WUxAUWY5au4KLJvA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=8112)
`pragma protect data_block
3l2m8UONmp/7H9fdVZbpxpmXcLOYUQ8E9OKnRpvBGbjpTk6ize2OafUZ5gNdSTAuLnqg5+TsfXqS
6U+Woc0//9zXRBrco5/eLgzG1rkrX11+hBKkW8wTLiwwJzw8NTEn3tcTZLiIhOB2JHi13Y4QxYXp
kF75YOr3yDM51YmoCwpJA+XaEnLUKXIXrzbMfO0e/8n4L3hVYB12Q0BkVeBAgzjEXmizZ/PfKWrz
mv/vKwlcxPaa2PMLUp73zQKhpfSk76d++ENWbsb5FITdK/6HKGWD9odmdEWjQEQwH3D0ufIlN7p4
xaPpaB5K4crzVNzVXNmRqJtqfX3/iteWN7hpPYCdcHTkpnsxjprvY7vx12G3zR/IGGLxFqmqH0SW
SpKzWUaOo5jyfnFVypOVgMm+lEqqCYUyGaQwY2MQrZwjcdk8cN74LnaaaNUKHHPePFig1k5AqqBl
ZciFKmeMnmL1vAPG6DA7SvGvG+3UJms+ZOirsvpa5M1vpZv3oa1xoFhb/amvHw9je7x0Gd83DgFj
BZXxr08cmTA2s9QOpZ/uwOxfjCKL+0MqvJj0sYJB9qXqf8yxyIn653xsn3Ra4k7bCPoAVTijUncN
bopx3ue9j4Rleke3/uaIYtD5BWkV9mUOit55WHFTtVZyvCznlBzpk5+DglJvhYDux8NYQGl8vbgV
UCh85x6ywrMqnZNbfF2RZi/KwfCml1k4ROwH7u/TkDVUJwkta7tzXM8Yf1c5SPaOrXza55Bh9xQP
myhX90scxmEOBWIdl+DRpXMQ++EaB5KDf9wjZBj1ZqmpeN1EOsgOuGupwNnsq6VLNY4wKlEErUYQ
l4aX7ICwuAXo9MyDYvdbN0vQir+vtkoae1QVsLRuhi63v8RC32MkNSVJ5nFY1i8e6ZJlP21PGQKd
P3oJ/RYZR8GkhcIqP1nkPBbPYHy/ZyAPZ0Sope8yYhJc/zS4bv7u2jZW119d/uvyd3kQSxVDV1D3
HgpXDtzKY4igHbPsRE9xp3ErBkJpPR0Xm1Yo3t6ZtGgT65+0qp/GOWTL6SLPl4rM4ckUxyVhL2a2
27FtZZMLBWO15v9oUwffAjdxy+vCmnTESAzZ1sXZ9DRW5HY9aNYKwWfgeXv8qWaIJvgyX62OuaOV
s5BmDf72DOOYnXEEDVWyJQT0xW8gG+JbpsZ7c7e92R4MEjGUFvvGLC8Wn+XA0UI6iJIgEEamJgnm
SLkjZ3ZxPEwJ3yQF63arP8tP+XP0TlbEp2Hd+B5dJVvs9Yu3s5Jk3glUiw2oSTOvWZjxBuDXSXfk
0ZdUZX5m7ecJ0dpQd3UfqK6+c2sw6FfVs3awU380X8TAcO5AGHj5dJGIkQnubwrEd/nqmVurxwvI
clE0MrxHB12LDwzdhxfCRwfU06hN003KfVoB7J25C2a/g+SnzwkOjOnxmrCIB+WQw6l2yO2oBakH
FbHmJBIoL0Ol5Z26SMiO98/B5RyTu3kLxkFqhUamUa9TOl7kHvPRqfld4JEvTIZO6/1S5hd0B6uw
7wp0FRNJfNB1tl8JQLLVGzskLT0eAoWFJjYCghBnhWFvyIZa19mCKyjTrn6NZGKdtlUPrFsbtF5u
+YdDI+v4l0+BN4CkeR4/5YTa50T6rxL2YAUEqnDOAqjpVGXM51t9aHP/GnXHuuK+SB4YJ9CTezqB
LUxpaMWQSxW4hmhzvguw+Dkv9daDtD7ntjhXi8pzZvLzLGaL94SXi6LpG56D6YLF80nxo+n7qRw4
yFynD7EaQ5p4EoilZ4scwQtphAatMwt7stGPc74I+/Yv7WNpC4RwKzmO8wlVe9gVq35PrLqDc0/N
L1zc9TSxJwRSAY9a3qvtOgO8G6RuTTc2nkIn0Dz0h5s3V4D6FK9caFefYLhv34Mm+2q/bf0RSL4H
SusqAv9ILVkAaodzXqvjuP9OjUs5e4ZSUXb8VCHqHQemNgM5ZcCQGUhvcVG4gP8DGOl29/Emi3Bs
1FiBMAa+ylMQE/Af5EckRP6e07if3pUFKkDym82EtGKGYkb6NGDIAem1GnXr8qmjckKikvDvXsrk
QYCnfSzNTAylZiiY8Mo9sQH3XRnuTcNhCKdxs8gL9fR4D6sSdAhCvPSyKvRS8zHCDJfgWOjH/VXJ
KMYwsTwnTSTBTmdQP5arOYBKktKR3oGGI04HOgq+3+oaN6PoH2bezxHx1LO4E2nbHQKc73fsgh+N
5styjqHnI1as9h/gRT3LQFllhz4hNphvIBrub7KlCZu0+eEqWAiMGZK34YbgjFQm2pD8/81Ub88b
UD9oAe4I5/jiSTljmRapJU7RtHNvkh8YLNyThcxCT0NzR5+v5KzBRegfKo7QLeaWVYkX725YeMZp
hAdStQ/LbkQzZHgRud+sW2xTyDpNoEc2aX02ctcM+fAizv/Tdm3FH2a1S3nx6hNGjEP6F8ZUCr7P
vgF48Tv1ZyfhTKbX/uh6rDB3ul6bqDFsrEJXfGKJl7UpouQoEsDhMXWisw5wchASoOZyLhUcGzBF
bzkXSeA+QjewWmJAT+D6RneX1McC2Kb5yuTz+FcJadpZU9vDAMbTPT9ixJ7eexlUORLi9OljzByR
AtD4XhLEpBVV7DLUZVBsZAtSGKiey0cfT0c1oFm1z+86gC/yRxfi7gWs7Rt/49isSJwvNPCb51B9
fGg8Lg6OClpQdjLDAPTsohE3mX91WWFA9avaio/mY8L3az+qHtXd4dNZQJlLCTHG5T27Xy9SWoNE
AhLxoBoe0I7y6wJ3KFgeF5+d1Yeh/MJyn7uuJ3ogBP5xo/gDuCqED4Gk4o91OIrGqYFXTHtlRckt
K0RlF8wGbO7GzkLmU4UMRuPmNsSYZPd0I2b8IeGYQyhkpsgCh2Ta5ArLzWMhLTXEfQzzhWD5kKxb
6EiCRpv2S+Cs4IABLECt3ud1XjPbsqneT5op3C8bB0Sq6Gd3f78oq///0ZbE95ucqSW0TDMuhH+M
JPUjlUGZ4MLAj3he3Exnpb1hTWoc8nCzIkj1lReWV9cR5FCC7t3VXTwMYY+cYQzlbfi6zfaDvGlO
5u4w+hEaDQxbQY3nJEZ6IvJvOxmO2Al46rvCqJreoEoQjuj3zTnMggDYcNkt1hDVbfQk3eFLZWCK
hdieTPjnR3HnjC+ZrIAw+5DLTxcs6kyz2h1DYeaB66S+Rmj1mCv6VNAEtar2mQ7nrCiaL+b0f4V0
7s4F0C/IRO/Wy2/Z5yZLrOEBiSclhZQMchXdqMqnpT5l7ISqaa39W4eg8YH1Y6Wq3+USp5pOGcpF
JohFqLPN0aUpbwYJQ9uyXgTysYE4axWyurPiRgQ8ZMWlWcLWRFeXE4crcKf0C/VntcBmoEL6hJ+L
Q8JY8dA1NYRn+KlI6nTODowBnCGkwn6a+YERZSakkPEdKxwKxAwzFR4ZOBLE1TUFoumWHnMHaHUK
YO5AerBVBgBEH3C4wymiwPLrJMiFdQ32a80xc0Jtrl4CIzVfbYYfGAWCWRJLUKqlrWsJ4QjPWeGp
JcbDiayMUV9SMmj912n3Jz+O+c26OZ1ZaT/FKOojtsYHp4suhMwfcqTe6PSuYafoIfKmk9X6pwd3
ClJx0zhbHdNWEjWs8BzW9OG5W9CHKuUedWQMfkF2JTDdVfFSYz+Adf8Lkj+HCzLXl2jdo8Nklnfq
4AjVLFg+L4C925+qqCdNMSgtBy+lanNw20cvXBEWlSaK3BEwAJHU67CkP2jjMJxurcwKtGQ7PLDU
4xpClKduKS5vGBC3pJ8aQ1DNS+khl8VH0ZBNQbxyfKTMmBwUXyZnUanT0HWQVZMZcjEO2illHQAB
aw7wtAtn1Z3RokkdGidb35W1DvXOcMcxS2jR5tEPj7qo6HenDgDVF6UFXUyx2fOUK8ii4BFZujQE
MBWaeXuyjiz6w6SvDaJ0beIMCMfCTy9ITctZwHl/U+Rm/adj95OQNsUYFVTgTkYq/qwV9m6KAMuM
qHcnvWDO5fBEPxrmFqXCShi+loAMj1PF7F/M8D5le95lO/ztXvjBMY+BJKIoOaDutazy80E0s3cx
J0L+a+2FB8zc8N6Rl4msFMwgcsJUu6aiFkV8Qi43lWKDXBm20j3zKHpaGj0Zmwj8YRwYsKSmeizt
t0slQ28KGcNH/e/UyzNy9XkZXeTKaSmQjozFWWgwZ8n0AHwrr7fsPSi08rxNF6QyILz5RMLYUTbf
L2xhL6jxFviSlBVOFnn0lng6hGBnPqV4DnjJ1T0nXrs+LB8RCS7/m8tCMi2bNVgqfC/nMC4NUOnc
7wDWQCpA1xbpgkzRGJ7F9bVTYDBib2FQX99OEOf+XDfZBO/j2z1HrzOxiwCpW17nlZBnRmX0V/Hc
WC7z3mik1bFjyTuojRohtrH+AFpoUra/q7FVGHYRi5dD+pjrO1IUVrkrINd+a4SfNPC6C6myUaNf
IzYzU8AMjDsoWOWcopL7yJqO5z1Gncd80V3vbOEDAing+8exw9kQcZIIuM/gEfWkMXqCxBP3VBHm
W8bTL/9Id+8zpQEKpRtBiJdA96xvaJknyAwk0j0Pvb/g/TrUkQzr54ZW4lGkPcqdkg6SAogoReQT
SytOvj7zOSuizaLTOEMfCrTcCsCLuMTYNUaMZTg5JxNFG2k5teFa4gB/y+L9KIhB3/c4xShi5/Dw
MPFhmgkineBHXJmyKvtY/9Y4UMeuDFTq7hbROZOwZ5oHoxUpskEITGRuHS70JjuZCj1oG6eYPhld
Wvz82cltaz8uHzE1uD+v636ug56fa40m+LBWrqLSx/8XtaHKbruKapcHgj97hPBKlMDwPqjoR+gT
Jg+upv3fwAnTGFYYlOO0jCvc7vxdFdXotB5bEsUYehpLYXFiqSQ3cXF5TSnowXJWg3FrZSzDD2hz
ZqiHAh02MQp0mpWw8C61OyrusCLBtre/hQ/pN8GtwPhGNfO2V0XbkwaeJo420Q8WpS/31AEgFB7b
mgdLvDqpINZij4WFFaoXTU0II7lJ8higAeDqW3lomtsVhHAJDfYVUUgWZFBttcy60i1j34goZUyg
wGn6DLAYORuMoT6umt4EVYeGZxg4LWwy9qK0m6R5HU5WZ+K3c/WkEQquYiezuAuBplVdTMHCG5u4
jqSRjVgEcICN84Pv0iJT7qJ9KlNlEnKKTXqnEhNJ2+K9zMNpevvCqjm5zu8Wz0zJYJVCGWl5hnUq
xe+BL0ecEcEG5zszZRY4GFEHyYpmvIIlJI2RwWcAQcQtptfrIdwUvEqgwELc9Al0G9GNljQnCUQp
Kas9K6IzSSHAaBmi290lUXb0Ah7fPIY9q9ShkyuZWG4bFKNQgn76ZoYun8uPYS/Mg2jGe1e6OHIu
XtqNGIA1jPnsvW6K5xVzwb1HOjdqqwOuYLqyvosQ17Bv9ewR6QRZpfpkuXCLEGGrc0oeLSoeyzaO
u3veLsPtkAzYZ2UVHWMeOzGwQ+AlPg3PU6BvEo4NI3Rq+xM/dDBxgJAyyxaJCB98efGqwleyDU69
IaFrQGtVIhJe6SWBTsI/t6LyFsfEu5mfnUr3wHaeyeFTjHhsXsK8wQcFEq3DTwlLRq4prHmFprxK
N5E3wW+GX6DVgq2VvpyTfkMNKaXnKutWO2tI93Cka/e4ed+0fBO32pYq4c/Sd0af4OGhBzED4OD5
bAA0pgiJ+ZAO03Jpqws3uh4NazQ0+A6MVJbLylPOfpvX9zJdzmFusLFL6nXqnQVLiRAgY1djIDlO
0ecF3zvg0J71qZucLA2EftmxbDzHpwUbRQJvzmenCtUIY1xSZ0QKtjWKJd6yWyJs6SdJUOqn5+FI
/GJaFkaDh79nN00f4/Gvp+vj7kY3z6xawUZf7xeUmxEPOBd9hjkhV5H6fVNZJ8snaukdOVMkF7vl
VWGD5Gh3/zyAmeYI4ONw53Vy3Qjn9FZDxc6j6r/VLDGLNo8ZW5vDWj6pBUIf++Vzrybg5ZNUpcr5
C2dneHjWSM0Da9fRdKI3NAh2AV0dzBH1/HJdmWOUKvAuS+N4+iEVL3yAxbMtfm+M1KhXLiJpWcMg
zP6xYu9uUcG7mi/ni3gHGWyKy5LB4INFxfIOmTpINTdDn8JfttbJsS22J8uOyMd1T0INKjtMBYeq
34253of3igUciSzw6AO9wNvCMw4PRawECBQwJxwmP411lCCXx99NLDGo8gMZkvGa/mKWs0sgh84l
7/4RagA1IOdXsuCRhe33YdjEw5wSNZgDohuwMqZd9OwYZCo2BtRONXSdqaYqclvyIz3NB+7nUxpo
shuXwYkAcUstq8HIgvOJb4Gwb/h+m1V47tyDZAppDC6MpehMbtn3datChc1ZASzVRjlmJ9dl9bYV
uGSRMEaH/6M4vDMxn0yGS1/PVjANrquBG25BbMhrSFfgXTyzIuwMezH20oxYFvzl6xQzHaiEiEF8
fVN8OX5w05woyKu5S3r0i0PwaKwNl+F4GuVlp2R4IvJJQnd5tIyC5shUVzIsIVgH+3dP4ZTjhSiv
gElTJG/FVHyrFwstUGfIdnXAtlkN22TvoXOuuNz2jWbCUMdirFYOYXMIze8b3Jrf/L59Z8AYrk2E
PO3HfJ+gLjtY84W2VMjNDdSPGg6lKFTXUo/wxelnhU7WAxRS67y1Hg+XEmrGHcbOflRf+NnFGY9W
ohC19TFrRcFpvz3H62/0EBlfj0nwYhIsZGYF6iSN6EiYwhZntBbc70WIMXqmjfMQeJZiciu3mRBZ
ZDRUWXsJTnWMR53fBdnUz+km6BD12UJngLC1VFKLlm0JJ1PZHYryfq7xJAFqC8cz2O7p3aCxTkLQ
vn4JrIrBmEICFtjhGjSn9nSs8B+2lBcWSmqnjNTmcN7gOmPsN9Rzj21LIG1Gt9gvQ0HdVQgUUNxa
+UlRqyIys5dnsPqpikAjnaQXu8J4kWdx3Z2zoI5ZX6/HZxon8jqwi9d3SRP7pdMpIKVlnkaZ3Wn2
ImqfltRQ5COyXV4FHI+s7nVCc7b2rRvQOBPPLGFlzflS9hvJ+Fe6axKwoauPDG0G9GENzR2OBode
yhmwFvXb/fn6X1rBWbpk9ooQAsy6ZC1V+SIVq8L69IXJR6zYbd60KJvPFv0HyYkVMsrqvw9aPuVj
vJCw81Ir3g5Xdy20TLDSduyWRPSM4mp3OduJru7K6cWVBov53U1mSQ2uxcEj29WA31vl20kZKp3k
yt15T2CwfpuL/9MzUJo6mNYh1aLCr5NXeuPcjX5xrDJRohoHb1kQBSd7QG/3gmrpuY80yHrdiHjH
uTrMsH+glNivqXilFqK5FmgVaJQ8m2JIVVOsULUVD59SqhPR5IvBOwpuqVXPA+UCr2x2aTiOaIzs
5EG0JYpCiX+/0bJ6Vag1LA8t1p8ADHvdFlmohlr9fINwCnKQ9SA0YxKgTYisaQ4CykExuSFWlOmv
CfP8ziKbzhWgkpmYPtyzz5wDMk8Wi2MA4zDS1fhTC2gW77W8JQvMSWTmu/D5doB2rChpmBa2HnBw
yXPG6HJB4d4+c0Xcvd2ZJ61dxuBRAedSxm+ub65qZdL4veBwdSbnQ2LgW/lIvIoV9prfHTL+1cg/
YbEHkz4K9UNTZxhfo7SIbSMKAT2u7MFKLSxXWFAH6G9adxWfG2Dt5YK4r2bBYe0xfIgHc0gMe2zC
4CsXMP7XuaQUh7sdC1KVCb7JDf8O8qtUXHTRFjsmJyaSU0GpoFPubWLhJgRrt0lkBZgiUPyS+oZN
5wVgSfntTHB1qzmYFIi3jvCZ2VQlXOdeqLb6vludNxdQa8PdY9QlbfqB97bjH2Q7CK+x1uT9pb5a
PufMHnaMk7EnGtnhTXcUpcxa+DOn1RnDRWtuNF98oUXPM1zAJEDWLZVmhlBQVCcCIX5YpioEeGg1
7wvbQLUTHsQonewggXBMwf4iaLRvpym4TOy2glkXMZkbxtXMQA5+mXQ9cRGewrfaOdZw7aRRL1DE
TmNhfACkVkE6fefgE/yI9s4aQogCqzzbJbk7zcz7cYVa0MVObyXOQ1Iy54fmUBAwH7RAsgR2k2pe
yBoEZztB7yqm9FjvC3ZlzZz61LVMhA06NbnMbKTd4YBzsDlaWCIJb2fL3DWMYVqvrHAyYHPhMIKv
SGQ228W43Wei2OmEuhZz/2RjZj3kPy/dpk5pWHEQleHR/SnZ8agmt7cNJXD3MkS1CL4Dae7iQHAm
kA3SdyJr/s2GNZm7F4IATFwjkD2ZJd1shxTkcL0L121NwVlNwJvDF0efLXKHb6C8SweFeNrX5hH2
Y2kQCAbDjd6Xj3yNeNo/hDcG4vaMXpjGvm06S1HRCrX1XNlSA623wlWd6LjhWEuXMtMKr0QiJ/B0
i2TtY87aA1BcN1IM+8BuPJFwyQGpqtBH61RHMzlQo7twFm9J2CyLafuYJiy8fGxq65QoCyAeZLJF
oAZCkkFumdnxyyVbg279L1PJ8kl8Bhv4xrF/v3o7GFvJaVItaC86xKeXo08HR5mgFy9DR1RExNJZ
q5GcYdSYOSOql2cmF2WIIrQK2t7x5Jcf9z2TzyO9CWEJJKT1StHCsfx+a4us4H+y6nS/IrKT3ADe
E6jLlGVPtQMtNaB5LpMiyEBwqA5tdKLWFa+sQdXUfZPWkyA1IpGLewQCV6FYaYHj38N49i7hnZiU
Nw/RPoR8VAOCB3BlYibO7U354uq3q51tf9Kr/A8g4Tw/GZc5jGJ+jV9j1uY6WfFE2NoWswoHaCIz
VrjuSccbvojzAr7QFODphTOwq6k9FDTJKuJE8wkFNn82TDrzoflLt2fIeusYQjetCNYTAC2NrxrC
vLYE5TNdolE1CXt3ryJDSy98Okzx97fDIiv2QntXJHFPZBp5muWcf8Yk5SMukjZvy/7SZhQBH+dZ
4iEnaLRvQ1qXXJKNmbwUr69AuzvqRM2oS07mGWOVA0ilAFuEjYNGmB+FgUiKLynXcH3u4h/Da9Vy
hXhJCILplawqw+pkoUEEkQB19lTWFpsU8SPbXXVpceUqitLftEtq0AQm2xpR5xStn3XUGwo1H687
3y7sqgwk4XYPUCge4Jj3Yr8N54anBFI7ihnLyDeDIpsVt91OrFkdF/4Zn1ec90CBkjKpWATaHHVX
/xj01OUPwW4SY3YHnk89r3uCAhr7RHEqHy4rjqq96fusEiI1bJ+d/xXc7xvBA8U2VmrLGQAjdsC1
7Uefl2u4cOcINRJNN5zDrkFvMpYxX6ow8kCSrYDmMxeRJdG091hxtj5l4QTFfqDjFqnaX7inctFM
uE2wv3Vit3qLyYrT+h0DgHp17nOyVH7Ci/eBMRQutWG/I875QM4k2Ret2QlpeS0gneT5vQHBcmIK
2WujJk4To4dTxYNtw20cM0bS/WmGVLAJ0Czp4A0ONCV/+YyV+O6EdGMyaj1Qcs3KXm1oNLyvY0J5
0lv2baT4ohkIiH9QvX5RxK1MD1ZoN8dR5mh7ejKHekwJOuERN9JyDG8lOctJYcZbUGbWxTp3Jr9g
DONvFBnXDG0YN0FbF46Dvy+ah72LbwCc09/HXVqStyWwvdmRfw7tSBTw/DB/eU+uaNKXR+1oBnYV
XHUf0H4O48Hm9rfVdSO1rdUSiLE73Q9dTJ/tXxCso+j10QLDXsPgmZizRsKaK2SAdLqKsNMyxtM6
Uf3YJ3TvmN++4HA3cCycQ4gsToYrcdPlf4IXO/UlSuZ9xbo8+2j9Ggg8BbnV9Cf7O9wKlHW40xmk
Bt7++tpAN2zNqCI7xcSymGZuHOJHu9MPi5r2DGl36ZQOkDsz8XvBGN7UbNpeenVDNAik7h6scgDy
5pSlcAzQcjQTcC2uhL1yI7heHovpNc3pYhWkh3+4+p0WgWHeoDUE0zJLJzKj/90EqCeq0CwdIeBE
tj9NyA5UpRJoKFhY4vMmpMKarB3FOKonwMkYh24zi2CJO71l80JDyqcDVVqiSXsYnHgVvA9yVVJX
VBmSkBibO2ArKU1Y28xAkmJbLrf5IvejaBP7Z1oS/oL83bMhP/z1lPneXtrL8KbQvH79kmk019I6
n0CHpANtHbbzrLglX9wrkiPmJBReVBoaxcY9HQIJFK/GtMaIp11TcuGiCsA4y8as2YC+nHpk1OOK
GUcEKFfFEhbLZm7sOvLlFHzruJLOHuGGaau5RzKhNarlq7fPe6OfA9DMfcUuYFuADCrF8nA+JM7L
3jx2Bu8iJSEfrY++9HVKgKJcs11Pj6DcWPr3QrHRg2ONENu4wUUsO6/fNiCdiwGrrav767oJHhDV
ZUuEJtFmpmiwrEBuML3dGnAY+S07/burMFMZW5JL5vZUZe9lyDIAcK8gydZDAFqAcuVi4AXpSea+
XdWQ3nn5HExhFC+GEZd0Vj48ojQG0g5RmLgbkplYFea5qsK8xV1LBRV5JlPz5QakNZC9+nGnNLfZ
wTANzMHX/iuMbf1c4YFmjPDw0O1jUu3p7xkc73o/Z4tY+OAocXKMlWv1YY65oFnZpcYW0CAIuRO3
HnWSkgbrRzjBp/DdK85WYGv1YpSJE11X/I2hN/FcvYuKTh3+Yzeelu6hzcqeZzUauIl0c3hTijJn
vj8b1X3dCRqcjAatu7hWCGLCdmEaum0h4DTnc+DN3oSObR+Ygha7chEAeNDIDsivEFKg+kMTfccF
iuQ6IPmxXtD3tvm/k9BeE6Ma246R+srDb40/ofFlGPLQsaEqApCQvm7e8xdtOZGF3OYOA6scLlDn
8SlerYVPerR5abUsxAIA6HE4HBexF1dZcB7MIve+ByUKhNt4nMQhlkzVG4RpSG9tIWGeHUlknOo0
ch/vA5Lau8wEEUUZ0tkzPc6fTyplsTtqlgh+KY1ZnwU/TvhRfq2BbZ9tPxw+Xa9jwzt5b6u627r0
hhKsLQOOuqwSkyuHe6lyIxjH
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
ga7z3iGMhGhga7TzPGleypVOHJn9S7KEP16RJ6j/y4QGRddc7/SJdXJ2zPvm8FTCqWlJhu6/s34X
gPP3kw7dN1YdiZ3wZ0Vzt8uhC/B62KTkMGylsJT3Hm/4AVsby+VuOus10FHgOgp78G6FqJDW2hD4
FEF7AvpJ8kF9S1ZR/yBaB9R5/vEzgMTG6H0b1hzTpBGPyaW1S33KG60mDs4uY1wSc9WkIOuDsX13
gE5v3E3AdV0s35W8mk90srPFan8A4v9WhQvKv0pRdTPwajKYNoHYw9l0a0ijfdCCo0SwbSJr+KOr
7KJQNnQdeGn2Y8dg3BGFPO1H0k02bZuSqUQ8rQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
dBwrqXpaPIvc4b2fzIcAYNKycDBKm/hw0N9OirP+O5J0w47WHpIJLrz+YZdtlXZ+W2OT1CCdKga8
l9q6LpHNXfMJe0tSBaUQJS9kx12QCBYd7pz6Zz4XteULmwejqAW/r/1SNtjKdsFfgoOhPbvsYv0n
RR9WE79+rnvNSo03sWloLz3If8EsTQUj+4AuHA6W5eeLCFFrjEJDELred9ftNf+GjbKQ4DD9VT1l
GYpqKI157tMW7VzaYctB1tIYsZm6N1scQY5/pen6aJE9XG/GVJc/lUhiKfjKkAB4R0V1b6xO6o/L
Z0CvpttfY2ekIVc0VuCKq5gMTfn8BkW7RjZNRA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=9104)
`pragma protect data_block
3MLlIGXYAu+SNVZUrN9axPWxB76fSavWP25CyQigoZQ3T579rH2tX4mOroKAFnY6MCrE4zy5SoFT
o9pFhWobhy1JNncmCcy/a0fRL9ZlIyjwjHAt323ZL0R5G1zw5cvTmFWPoZX0yo775l85Oj07XBYY
i+0FcCRCKdgsQGwhMUnpc6ET4ttBmjQUuxB6g1Afy5ISJRNYs77D5E8aOFrmzUzDFsE9BGcX8wUT
bT4zFmjkBZBQ+KrbdhaUiVbninMVuzKJe0egFOCGcc6CdMPwZP2SxWGkscRsjPCAUdXGIydg5Z31
50m/zUoKITRK4jViYvnHt4f6sELIUTWEwPvxSg4M+j+wpDH8hMQC98bpm495w9Lz7AbFBmLBe5IG
17+sbfU7k0MY2fUrDvsniZvkyXNkbKvNrkm2E9MAmf3uKtqsnMU/tF2um9tYyMuoXrnv+cf1WHME
rcGa/NDEnGr3zL8P+jWgeThli88TgswwgsRldtZSZHdEDO1R1Eb97kPR2KAaazYlo2Q2STr+5F6V
SY1q0ie4TtY/nmeVptSZJNGauW3hhgmAK4fuCh0LfgbkBsnHNuCX8t9sRAwVUkoEOlvg+hIeL3ch
IbMuCTBsi9ym1EZ2NwdIt6YMzhAa6xgt6mL0uQSzppyrK9CSimYyzPbah+kviBaNcZ+XJClYLFwg
Dt034rBFaffea3MI9/T6EckVHZwmBgwvpnfxe5dIdxVZcMCrn14d+8gHoeJtodrk7RCejHv+C9Jn
yRjIaiu6w3mbAeAL4r66PbCB+S92jMdnwdBtSBcwI+pRfl8Y1ZjnMUax1D4+e4G/2vS04zWOHJPK
TAm5M/l7TRLujzCl4M5tq+MN/Sl/TrmT6Z4/ZBXtoFpOHicvprtU+bB6bA/TDiQ+wyauUCUWMDnD
F2sWssLTcUSqWyGH8nZQJkJU1GRznsjpDp4OUZFEoGr1SIfqUXOeUdRWE7kTsTGtuLLkFRULD9ZC
icKwOzgQXLWvy1haIHsyX6SZ+d2z16A+qjc4h9yGuTAjU8NLa0V/nk/gnsMB1qd073hph6QLxLJK
r4sFXdYNYgCk5RaS44kcalofpqStJQULijgevhq0IIAiHku9ZgDSCzWAw3Mr5M2bNizLX2XXA2zw
yD5SKKgh8NLJ62Z1MJq1d/+XEurLezROXf2MzGpmtx5eT+YNTMToyw4wlcI7tOteLNTVwpN45tUQ
B+wyQRROLfJbya1slSCz3CBx0TkfIQfh2iiO78hl2uIlnw7hygM5cDhSSbRATA0xa7ahqhvOPN7M
cHlx2JtFdxdsqSaZD9QoJ639DDyU3Hou+ECwMn0csUSwgAS8rtGVdP0Of14CplgwrGPXstO6akKA
3u+imfQ/w8L/PLKXBmZ4JDbURy7k1H6RKbw37csxd/ZvrS/pSmIkcNCzp/c2DuOoQ7gmrvF/T6P6
o66nwV4BSbtkXVm1Gd6pj8kuzFas4d8qUgIJYtO74n7f/EHBC4KRyKr547xiGiwhk9b9qd0mjPKY
rhYsYy9gXuZh3r68RGneNEq01MvW6g9QFwK1ZOIvZDYOR4QWzSf3jaria7TfeR04B0hTDmN2pnIe
G0GNQyny7szBaDLk+3oC5dKi2x7IBMiFePNumBGpRQwF3BZOBafJAtsThr6J0+IuaIyGTu6q0CRE
pK6/stbZUIyDHLZTtsEiDvCUoqJt1Nwycg1jZabyqczbNym1H0NA+utNZBXESxVE+E0tL5xp64UF
6UUd+qxyLwKovERkzivDR8GuW1zTirEOV5S4VxepjAekJHQRl/DLLebsO05p1WmBlr64t8l3I2Z4
eBoTyoAckywhyY3Hef2UK2jwBO8dnRLD1Fu46o95g5M70RM/CdS1OdLKSF5ccJEDtzouHFkJV1Uj
jF3ui454vNAg2ROOQ3kKuyo5BsEY2EVCu3TpZq4c/q9GQLsRGPOnx3VcTR+6BZb9QBmDwr5qk+/F
Mfy0nKqqzp3OK73AWybRMjmJczTm6ffP4zxEkfUdzR127EO+OljvRItBn8LSuKgqUpIu2NxDCg+f
A8xmKgcdP5Vj8cz+tus1NipaLcnS3rd6rslS/DaabQM/fOpx4ERbftZUSiDhPxRfGlVjhYH1zMEk
pr486KmY6LfVGaqc2pCdgIkuSoohsNiPN8xmmK5O9HjxRm7IYdaUIvotow0YeYsJys+80/gJB5s6
cE/ss5YkBWNMAqtri10qAqP/lHRchjbTFTFInn1auRmyFcN5WTjU9MqXhbmBIpJrVs6hQ8bjrGbe
udyynSp5mkE0eE/e2v5I1wi1YhxlXU/wpSQkq7AW/DgOKirxvaKomORblPuNuqND5ETjQo+jpEPM
80/aOZIyPqN0aWmrTJE0jsjxS1AJ4MOENCzTG523Wq1bgye8XzrN4fo53VpdHD6EPKSh7ZgGV7sq
giQ8mzKHA5CetG2XXI6zrPk7Oe4z8m90oe+OF3HP34C4sTOp/x3Y+GqefIC7NoHPNtvs6PK4n21W
QJDfypWh5VF59VtNEgflzAT2wYDVtih7VEgDNBwrj5ychDhaeRx4+0dTJ9BZTa/Q0qZqOY4erpsq
jvneKxGNPh7zRngog7RWOBuH1Hi9ahuIiY+gEC8RxoTw0q9WCloHfF6cK42Bey41W7Nkg8Ic3W6O
AV81HlRcI218/r7yKU/7urKe8KAq0lmfWI0uIobow6NRr57vlBBhnMIl/DXynMAD0MicHsH1Dhyn
h+XWBoQuDUWkaHIh4zZ/+1qRMEs0NnSiSUJpOxoccGc+tyhoKIypXhHvUevk4IqtTmdXqAG9BJVV
k5OY9fhhlE2OW/ibdkZv1N8TAqzbACTxaJsG4yd9IXNrWQH3memdIJYipNklf5EjC/KvbTm5tyl+
BLxlplNCoR4T5q2klsjPNTl8nKAiMYCZJ29rISm9ghJjvtpxxC7iQxNuwy8DpjfL8Uf4MMBxii/H
GSJtEZy1R7DGqeOvCIAWAjS1+kkxdMrlh0x3ruEo2+mWagYuF7zcRwv3TrcxsdpZpxjAK3KuJQ5d
X94lkof9p94Q9FjBqgLyhEjFTPbeSIdMHrEiuPoqCq/SHstw6UAe/HyD6+3m2O2WR1U2m9uPatvm
sJxRvmVVaHWurvpn1JNRY5/mpZqXlkjzuf/rk4eL7YaveH1F0WX+Ql3Pd0MA4RpPOCPoYJ6ooi3X
oVoBCaBgNLwuE9nJoaTWldtbdFa4ZaDZk7rQMlAKVWXu5XPEChTjxfzXr9iZw8Qdf1rTNBPLxMWO
LS48BLsmr5GXjy67UEUXHgGbVRrUX2AYtWS9hX1O9CEOcvgQiFyWG7+HS9TBB6SQ2461BLLzDSIm
tHQ82QNlJVtLqGTo0WcNrWtZBNk8qWHaU3vXA5QOlhzZmHw9E/y6jLn511lV/OUgJnhM+VkJUv5u
1GWSh+SGQ7IGzBlp1mAMXXSKsY9cSzVqiU7ytCkCfz7j3DJH5ntdAicnI7krHr+QdHoHVl3cPRNN
NTik7Oj2TIhkPWTVsDBGPqiRH32Jtk27wkbWFHmGcDeGjORj2X6SeD3i8lDS8+Nyx002zkXneNjl
oDd24LPJJCMQRDT8cPvqruaCPj5QFhcMM03UDgcEe0uSRvG3XOUcYyRtYIWKz0P0dGmT2z7cqLW1
ENc2s1dNM7+/NGNv9+l1i4k3SUF2wgInwkta1RWKB56XoibR8jb9nZfyKAZd+ByhormXeFYgJY6t
2znXbQtUxE20pMTeUchfKGOWsK9utDo4dH9Z4WRPjSETi5BQ9WSSc0bQPgwEkOS8CdxdbDClxAUe
3HXKO46hwViJSBPFmhQVlUuSkfc/Qx/KhZoxrEyYemgMqJtdSQnbk9I9GnaIoeDy2yg6S2XpX+7B
z9BB2oh1S+xi4F9PofyGtTO3tcBJ1/Lnqflfd2P9J7PrJ6+ZIiLxiP3RdiZ8qBl9VsKEPgYsP6Eg
GVXPNHLc/YQXcak7ugFdBOg1QHcWgXJ4VVCEvtoDFFzAyqlHNJ12e2cRpKFTUw+mmYuKKE2X0liZ
gE6AgMehTghpxhW2ZtNCsUDiE+XxzmFAuXwR01pH0OmpfYM5Gs5+ql0zq2OiUXv4uAXgJODLW3Oo
UMp8LNmKSgxn05S/gvg+CQv6xwIBotAlitUERe/scua6P02LRJYK7skFOkC0gUrUEzVoQkeiXqDn
+0B0nQ5+lH1aE580e/0yq961UMv0RrPJ62q+EbmZyZwu5ixNORWQjC28sDhpEBVKzQbyKlsTl3PR
8B5px6/m0sZqtDFsZ5S+pWITdhyIqPvHzfWZsomTTsHDA6c0l5HDL9GiBFI0HY99wEiKzOypIT83
FOxEI0HugnMVoH325uESJ0tgly6Vg6gvVaegAdfYZYnWD4cUJa/YCLI2SolgSSY6/HUFQWZPlHSa
uwytlojK6jIAi4ZTJVbMCfPCl/ftu9iMtk7QpMPCbJJ4+3Y4AToXQzG+F5En14E1xcqTz8QeAz5k
MaG+CLBnoBIeKAeYw3om/6KzHoJT4qAzUhO3XgIBkgHI1IC8PzwX5mDhqVSfXEHnKVuwleq7gziT
PKscWaZc2Xx0KoVvEz6xdNM/GTu8l+cz02Kuz+vvIWmRp5Yk6nBt5ZdX7mfvPucGxudayGSNyz4R
vTp1wdX+4v9BJyWhn84CMCmj23gGuyl/h+hfHuFP3rDt3VlJiYGLRrYKpHxrSU6V4FF8+QfSW47P
lU4miXdAmuTgbQBl/gUZnL4Ea8Y8GJd8ZnC7vTFB4+TcBhFOS57rzr6vcgOwksjHuvpnSe0+v5up
/qpQ0BUiDjXFE9ioy5jKZvlAPwy877pIuXSF0s5Io7V9+0Gvj5ywLtj9om5Xa1cc9IRlkFGu8VTo
gloNpftvTYiLcgQ9XCkRez4VkhK9OeTUu7hcF9feSsIOcPxTj5nup38GVnq+18FQXm9PWgY9Zvp8
UKIq+ZOt9jK5lFIg3PDPjB/H0YE8NtFYtJOYTOCpub2VQtpl31pdiLRMMtJgbVIhVvcIDSvLrK4A
UQsWbOKt9kK8HKXchbzKQE8dfnZpxFjFfsxt40CT3oX5g9kpOfb+hLmp9OPjA7yUU0OLssJ2BDN+
lJgtdgtPc+nMgC7np7fTeiYz5v4y/cA06w7oMRFKgIIeNKvplnPD70X0sdvIieUSVy0VBUYrqb9f
AD6gXnK1b4JW3DzB+S5sn7P1QlrqpxgPsHyZA9QeY5fYRSW0omlCDh/DMAwKAf7BJum1e4ToZAfe
8pfdpqQQDN+KIEpZ9ljHZyN++7cj4D0MmDQq2eCYgAdbedXxAQ0nyNK5GZQLt7DuU2iY4MXiV8Uf
7GmHl3w4E33gqnNvmOdqmVAEoZ6m7iN3Jg0Pan+AASxzx2kOJuU7T+GiSznzLMvS57lMvtN+A7iE
vUIXWpikdFmytaf1mGV7oi12xlmMP6ImwMvhmQ3uBSaHehqod9chaesceujXyFbvgaJiSuSMRpet
AKC+3OrxT/FcIZ1UYFYbhyhzf5SMuozNs6TNIy1oyuTjo3E38b2dca72hunn1ywT/RRHvgPBhxZ7
u2pWNBJvkPfQ67GvUOXnq6fBgUZQOKpQlnKUjHU9YqdouQwBYeE24DfZCe6ZYw+zEdmbZbgsgE0Q
koPILnoPxCm1zCzpTTJ87GF4UZjsBYp5qxCWKcWPBDHesYJRXINipAm3cLjTQB744dOIVr+TaRMN
qeZJDkU0XpYUefrh9qhDO+012nvYSNRf+k+D/Mk+/ueQptKoDdqBtDO/fH2Qmz4+9n5STqyc7sQN
RBQ6KcRXCINsNCAWgL7PrasmeIUfJ2fWObYI52hHHj91+JXbtNYeSJ90HQlfeWzb8o+sHBM3JL+9
oeQONGWw3iIu2duhADUs2yGzTpTi/emiiwFsIo9dnArRP9A+AaXdiaUMGhySnOVgOfpJpJ2i8fGF
73w0fTT+RE9GiXdO+8sy2hnDBbC+SKySV3Pvyxc0V48762+gaatZGtrWAeTnd1MH7iSEE4ppxVsA
qf7jYxK1osfF97bbtRRyYTXGgaBiyiHjC+OIz4JIb2jjQeBHvm14gmmDe+mOS1ACN9HHfztjkgRT
VvkuMx1Q4XH3naUMI68EgKzU//EEzmu6W5qkcKHYOm6LRgWno1RVkzyvqx+UW5cNYe3V2kmfn0nA
ZeGN97YrzUwxmJBbRQ78YQggdj4Z9hUg/abJwUqxqOse5T5tn+NUnX4PpBf3Emrqr9n4tYPMmq07
HbMRhAfFhOVk99ttQEWLK6eR/EdTpucr7TV0zTLUe2fdM1/x9IYeeXeOW7V4rKCN4jMaYPAIW9gl
VAQxO4j5PgYI+OHXFtOGsiQYat4kUEm9txb652oRW7QeSsjdxPL5VpXgG55Qf+gxNvigPhdKL1ia
2Gb4sDFnfbCCeW9Hs84BnCk1VM7yww6trr/HfHiUrONgTNof/0mDFuYXnMWG8YW5PV84dcStxNfx
JO/HLVBEUrL3R4ZNIQV+BMvEWDAgJ5o5NXEBpGlCYXPNtZvhtBvb+k1PK9Vgtwimv6FmnIcuwY4m
zMcTiMbDFy9oHSBd9CODtpqzuaj/XCBKoGVeMRunnoCqo1OMDU8QO08fIKc+R4IbkJqxnhn1n8jJ
5ODghW/hlzyatjovXVT0eMY+Bd3m0c1KWR94NvkflkhRjRWkH8KkIvtL90fzh5iyep2SS9jFV87x
Sm3nrAZWSR5yriLs8n5ecUn1R+FdCrGNNewxJI6i/V83zlQb5hjQOQyLE57Bz2d2kc+g2GeRn6mu
NSesncoOHHBXeQQQPovpR8apeYttoI4miubhDIKE8fhJHCkmgJ0nRsWNKkpC+Cb2B6sDKtC5kGv5
nxGpOVCRr9cb5W2SpJPuhr63LIQGM1+yef/b+xdkSGNDpIHGsC66MsOOII8pa0shJQL3AFLUX3Bn
l3rwR7LbtTb0r6hAFUsTfVdUu169PLgzR28bFEQghbA16YiWa9mTgyj1b/pFvL45fkhOIpSb8iHD
NxmhMs1Fcqe9STDqBnTvVw3tMgJfk8LO5wimgvkzctStRyTab/YzRChEca1cWPZL6AvHJWq3o3pZ
SDwgbuhVyIlB0kgwB9xAPtAW95FdNn94Wma6Yan40SPPot5z+8qKu0vQUDo+LOfsvX86EJupdo/F
UJ1HABbRf5wga0OmmYnL3AEbn7x+YiJh56oIYe1hzeqHutrf21hIRknge/oxqtg4KuV9T/l9RJT8
2I1mhhOeX1y2zDafrojZZeI3oAUaSckzRQn3K9OWJcwaFlzKgeT/0qjBLFB0Cd/N26+ty/nTrT8A
NgwLChezgsy7fOsykJ+hUKvNskGDBZmrifpGRw9UDDiG4H8bqFacK7QDrMsiVgMyJqJjjDzu7UMe
kn3YSe6423Wh4Oh7UAnvfaEnPR8xoQf3bHEsN2cggH1GwS5TZJ2J46W0pAHISc7vMgvIjOQU9U1p
Pe58ZvE+GVraKmR1bgUORyZnlRo5kB5SHavl4LD/uKghzV/fJbgdbvyqest86QfvQYx2l15q6GQ5
s2teasM9aAAhA+FP71tUAb5bpyDXnVmkeiYrAzDJnvAVyzPj/WUHMu9Ev8A/w0wyLHvYPUrSZ5Hg
s9F5QInp6gQVsfAKbKk4q9S9i2L3qD7tJSnpkE1SamAs+WqbOKNA6KHJkCcWpb2n5BSgEuqLT4RZ
GJQ3KEYu+rTvuy29gms7P0rLSQ1Bij5MComeLR1BV3mB5AQakvWi0FanzTDqaH6QEsFV7oTOAMYB
qvFqCuC9ScsIp0nugy6sog9jQ5RpL6GgeIlbRpB1HY965yHKrJuAZofZU4bpKP1dLIn9k6AZyJBS
FqdgnJCsNPURMwQnhFMRweqK7aqEus5RHmm3iwrR7qok+UM//+UMLwtSbyl5WRJ3u4MFaFJe0Fzw
biCRdbbmIqz++7msSCEsBC+Wezf4XDayQA5OPCBhL6brG1Md3AV3B6IMvwbIMVq43NEZFgfgZGbq
P0qv8aYTTJaV/Z+UkVMkMFJ/WFd0GJuZy30jgLh42DDDGRxAjBBOh4zTgvSWVMQdgV/Uiig/xH7m
ayxu6KAnGJN8k4v2zUMRB+ApzyHdBrs4OxeWRb+j+Na4E7xwMHy7XqbCRhSIz5biFs5ySpldWo+L
HDuYj8RROjLcxhzM8GSZ5nM4z+6Q4us953eCaNZi2dJfq0EAeye0Zcpe7+ImCwG3t1UlhvDVlYew
M3qqeu71H7BPZDdBvoCEgaEQLKZrAo8UxKz7lLopTRbNLYXkMupvXU9ykfAlMW0REaB/hwBfeuz+
JJ3aEgR1bhSEtrVXoYl6dyuYbGmMksmx/UX3Soj34zTnnTJ+hwH/IwgVPjziMAmbHLp2okIhD4k4
uMww2sGID/AvUpkhn8lFF+uFbslLmfZ6mElOJbIyqvx8q6x56hcAMAtuUBak2yo77UTaWIQmasWs
cggXHuPiBsSZeB8Psh8zfWMalZs0K4XPRqB8WDXmMNTjVDsoByBW0ulJvqiV7VLks0lPBEEqu0wl
H3Jqt+7cVQq7kdQ0IPiG429YtGIZm1s/UMZ2jG1EyUOJbmT1PHibm0Eu52uxM0g+k5wvTUrRXgVE
D3tXxdAiHekCdEI3IYB4qRCxLY43iojBpuW9weYI474JZmxP7h3ELD3KCtPWP8ZU8OaI3a1/g7CF
hvhid23xXtQi9dz1cyeI5Eq0vzACNJnjomED/J/LeBX6ySNfpvhPI6aBgrNVTPEfEhiBHAlMu8s6
aoIOYeiiWBA4w6gxud/KZi7/CG7Ej+Swsp+aUavJkSDnshwFiGNeVevtFah7Q6pBdnwQ7SS0VP5H
Vb7ryTwcGU9Q/LNnIYCHyqGH5ARtnXRJX2lGMwf1srtUq6qT0ruw7Pju7YDHklVXDZctH3LihLwM
KBKGt3cPiBSAkWMNGoFEohNF2vHOYF/i4bfFGuKkAneskFT/9I1zMHLedz8hp9aqYn0X+/+ZK5Ep
mZLzdfMMNPq8x5N3Jsi/TvlONHtHvchWitdNBqYKwK3kiG3apu9ni1MXALcetRvQqQDo5Yqr1LPp
AC+rfeBDuhshFXQ9M3EmozggnrlvipVQsLem1swhkbL19LHd1HYmMfUUxKCvahxiDBgNmnxG5PUd
mV1VRFxWHyePXhkQKG/KWJn4IhmLJoGfVOn4wRaYZUeXE/YAj3OBSn8ZHFD0sQVoVwaLG5hKL5nA
JYEl7BGSSn5AYfy63SnPCrwfj2VTNK/mcD3xQyfociB5IqSytj+1uyOC5PlskTLanFzrPLTNVE0B
ZbMkPfukK2bN5jP5TluoaoeJxHIAjFwHMnirQ0YGYX43TasQ2sdWQd79+5V+5opSCdMZ9k8HFeEK
wqoUkdGJQ+VFEmAQMPDLKe71SvnTvmi0z8LKj9FdqhglwNzQ23/xWA0FciosFPsP2GYKMxrI5C5w
jXZ2AeCuHI333FfOfiVoHkxm+EDbVO78eZ6Fs57tAAjW6wjwyr7eah4OEpbt53hoebbMR6oxJiWL
pEL2iehBcoLSaZ21XofJ+haLaLt8cgCXCy1/62aMvZkLMmHxMF0omPg0eBWCi/RfANBSu896AZLL
jplbq3OUmShHULzXBD9NWDyiQAoUXir51/auJhIQY3c5nByrf3oMMq2LwN422t99fGys5MHQ4pE0
9Qx9VRO5G/+R+DGNaWCPhuR+9cvQYiD/nw9NGjAnMtUyj4ZYRJ7orLPSGr9BNnKu6mPaw9CUsOgO
zEcG8fAoz1zifV7ookX+2s+gVL76kzIZMUiNW2jf1UzFVMIcPSHmyOVM5A46KOZRgW81dO8a2Jsk
p6CKDMFD7pwyah2BUfZM5toD7EUvWlEAjLQlBJeIB1SLPoF0HQZBRaouoV3KivEvZMg6aOg2+FFy
uMeJ7wHpOkLDKLJeNhYWfBFG2LAoNcx2r8p827aqCu0pTwNB37+kGS9dTZUwt6f58OdkV/fnufq0
h5MdEyBiJSlqncxxUUtR/LmJV1KSevGo8RepWiaA+2CUWVe817lPoSnGbiXR8jIrq8wRy2qEVgu5
2KRKYwbnRULsUSlyvicEZQi9OkOqsBM7n731imcIEg4DL3C+jTPLmgF5B1wkhjLQHDvIZFpJFubi
YYtAgRlQWxWiLCjvSUTEP5Ub3Uk8WuLd8Gehu5m63UdiQuCdE6D/yJfx/+up4dRQEMtXD1OuidXS
4SAUEJuI72evrbnxnYzDh3Us150j6Jpal8pe9A+qs5oh7GC/HLHjZAKJwpa0tz0Q92e7bDp3gWr5
t9IafGE4pQUM6wiaRUAqv/pA4yOulUveX8jqyag/KOi/kXittHEOaV199Uykk5ZDfCE0hwTcFaIE
dslU/ahdYXurrHxilF8bEdNjF/7uU/HyK1ow4rXZD4kEHx/0TxVHPeIQY/a3WnZNVRw2JPa0Zvik
g9tZ5KjSaf0FFgyGwb9p9zuXDK+9mHL+1GDzg5auHK1psLQD09Q8gj+w66DXHS9JS7v7xwLfqxz7
vqUo52Z1WgceBI6tNVHSJ5GH3CBXcicUjn/9xVdRMePo50b+/bnT4wc+lwx0txkWyKBxts9aNNAB
aY03xJbkTq79j6zDyZlFTBT2wuLFXXLH9ywQ1CMC3hfDXNbwhbxaPHyqQaV0PjhaI7lJDqNLTujK
lEbmz7PrYVmxmVUG1FnZ9iEOdAgKWyoCS2jC0e7gj+hKK5k6MYvFnXTmGGtT18bk+kgMCGKtNe/3
8fnSU4TtZWlYzAHKEYPFc2BA4PU1AFKUPsAZnDer8BAMCJ9kcgtdIX+JurjUPTHpYjUD6P33WYg5
70JdRTE3urIZUe03WWGE8xT3tYXuzNd7c6dmvXlPd9coCs+cGtx65WBak8O4KwZHAGp2URby//WZ
Hv3GnJUtn0/X9qcD4lMIbEL0rtFidkbluZ+djsVbIotaCq8UcL/89VwWt+6IllIHJodwIpuBQhVg
7mhqKasGojCi4bplXyL8n019j61HbfVma4ITNRo4T59LqMSROzOTzGBwhyjKAbY9sFbKgsMH6x8T
vk0T2ZPJThwoM9Kqaq7SfkqrAGN4PfyT8Jo3/1xxqlkDFtoMlzhDc1eqKNaco/VAV5g00RFoznyJ
eXv+3GCvJ5bndbEilWE9c3TPzK2pUV2h6xxguYTdWTgaQPX+/+qhhGNrv4oBqg6Aihqx4ZltAt2B
2e1lQDgFc2BTHXq0VOOhFbqeEC+Yym1JGucXX0ScrlACRTAWeuinhCM4J5s7mqF1R1aQd5UN0TRu
SnWzUCAdessLPZ3DQLJkPRtipqYNt1J3GPZFZFVic61vOnxbAxtJhJyjQp2MYTHUy2C0pRRGI1Go
uuUfXbHBk/WCRQrDZE0sX4/4P9LwiIEjAWT4m+pjUvxmwIeFgF6x/fr0hvdMJ6QeLZ1PKWYopAj3
FHQ/FEPZP+up4+Etkl9MAegldzMpXBfNcUlT85tFEt57fa+P4CQuS32XwcAuADFoaeKzwD5ZNJgi
0sHb2fY6DNvemfpgBgWrAUXEKtLpkZyigAIY8weVlr4+mhrD9SQjxmWs1evjzEME9eCRl0fBzvJ/
/gBywkStnGu2tN7uceQ9Pf3BuhEvGSpIVhjGml0pzcRK2bkd0+FAh+O7Zen6aXJr2rad37EUHW6W
9bctTz/dbOvr7ri5bvHABZN6oInExB+rmPQvI//MobMLhhqRR9vCs7+dThDEbrWG6srFenM2AwOC
7qA9cFi8+aLEhWtQXyYa8T4MdtBQNjkT2H6I3Fxo4VQy8OzJMwrSBi+0ajvSQvYgbyVjM2kLGFHj
rBnS8mJHYSG2sFSVAykyqGPr/AQg0vDDe2DG8zy/Ll/1m/pnXYzC/CN0uDF0cCI9u5yUPKaNeXJW
ftPdQw9oLscbOMHX+e0FW6GWVdJVfq22+ZYAPzqwElRAiSxqA6f6nYm0U7Wz3viw1uSv1haM7etD
bu0QFEN+dtV4ycJTaRBf99yY2G1N/UkEfGq7yTZ7OjJDodU5RcorKG8RsKJEpnFVm+GYrkt3S2j+
Q9krFN7yIKrSNNwRlSiQgStiUj36vYejOryEX1vdh97IPuN/lOsZn6+KzTPhnmbCnoB2sasygwko
5kP6T1QQsz6xSGPWKDE4N2xJcKCVNQ4PxYcRXVkt+qSclQf0tuV4kSc=
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
FF92Y2BScS1tYCbOJ6nl/yrS9tO5nLdkcinIUmduQUlX/rEFHoa3Ivyk0aB+kXloe21LQE4kGkQ6
Q9+cOvbtZsLXojH8eCz5LSxZZmj1OY0HgImQvBdW/AXKvPSh/8qp2AkQS6z06aDmakr4JM27sgw4
e8FcV4tuRcqkGs7bb5nTeggXj+gCM8w1pZjupaF2huj2/7utBwg2caonPL9QnFqNhJnw1y8cEijm
U2tA1t1pCHmc/cfMmTL1KVw5knK/j+GUCQdryhHqwEoaWgcU/WsJ66DlhJyiBG8LqQzPrvznCBbb
LaJ3ZRAbBz91jljSVrMpulWLCnotPmY5QRPBNQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
cqAgpvQThUsKP1YQSQ4a4I/shkrWufEhsDBDReUcDIwQgy0J3zK8Xf8BMFoFrewCsS2KNDRzQ+ER
jCDGccgdbKH/8jqChdozG61idZWa0ns7506SogoQlXjlqxzJaYEQMyNxDX7Ycmqi2PkN9cXJyFzV
5txS0QofbL3mzPtdA044rsuP1fkQj0yHft0ysK4zktjTKWnJPMDoc1p9qdrOCvbt1ZBLB18dsflT
y4tm2j7ie4QPZbNefa8AuI4j7gxnCkSCkqJB+CSn4ks4ndlDn/a3c79q59d4UozEclqodJLD4obY
Qe0wLjtJvGaBIVSj8HG9RNO8kRI3GFa3bHt0Iw==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=35120)
`pragma protect data_block
GMWtVErQpQVB3QwSqSu3WLxWBruia83TiqFim1P5yomKZZiZ6hnfn3K0QDrmVwY7PiE5btr6uUCg
ASvl7Cy7cI8Zc2flo3CREyieGYWShD3jicsOWnhG9bJjvs/ESsC+6mByzLOMKaja+OOOyq2GcDl1
cY6TAnixjdclw2RuHFaiThePff/tUT79KvAd9WuEJyi/TU9blIqQCQL8YY+IuRrFpYaFcJ22R7+8
i/TffA/yqvmPlssbcuHxwd7Novy5J3eqctKvenGtBr97c9O5eEAztT+9yTanMO/ruuWLGDgztEiN
4/5tpmubkSmnlgPYLOETdvuf/6dARPXfmJWnPQa627x+muA2nU3Ei8/ipVJRuFGJysqGcAqzHGHq
ICMFsr4K20gdg8Ner2KmLtlaQdKKX2ilB3iWOYxDfJugL+B00R43cgiT9felfDOSgwV8N2MQa01X
wOidkZn9NIq2JNm9Gl2YMJCFrsFKNFWaN9daEyRUQt3m0IejTtehXQH6KOuoQ3dvcUftcx6se0Pt
3yFscgPK70X4o9S9hXus8uyimjv1SMPIMbKwlTmnwUXyaUw7Ksu4j76z3kX2DtALTvRfp2PQ3Lj7
OvHlv+iKg7oEvoMVrY93sbnbDt/2UZy9+l/L65Eb8pxMOAzrpGEuFZ+stow/QjqyQgbJDvdqNyW+
iSZUoYyShuxAG4ogbCfM3M2SO216kTNCgOKdDCdQRgmHtoy4rYxcz66OU2pYKZap+LEBlhr8Enzr
bSfPPa3+ApSHuRUE4c6P/i6zm6QVqT0zs4fNtsHrIqcbzfU5ldrnCuu0P63UW++9eduY4rhauVBb
nm2bzBEFgLkZpP6mgMlAdD9ALw/7Xr+7fzXQgO54KIn+Z0WpkfOAxXWjrJZw2+LhxgtG+o4CDFz4
sXUZmjuPK3QHoHGqM3mofbC6Jl7QHUf9knIQxZ2v5A6N+LEER8Q4KO+ywbVHGh96TJwFRPzX5o8W
pbdOWjJyBdgUAjDwbPOOodfz4r9nWyFQKKXfwPEhLSrcf+BcLXvJqApBJYRge//KoccAfLGb9XBG
FzFb9/b84g9kojyCAuv8Yy9Vn0U/OJxuASNhDUsK70vCPtIpR8sSn8KCiCsDKDFu3aCrpSoLRLoP
D7B+YQp0ZLBcfzQvrXUSTRRSf/C5PNeOAFFaFdMIZnZMXrI7VYfW4ZM0HfJdzmP6TohgFFwMLSnh
kT9Jvg7QOXHvp7aT0uWbjM8kfC8gC1ztAOWkRGVR/faxnkuPrac5LQJUGrvbetUCVIK+uxrak8/L
qXKXlRdQSjGDFy3+IQ8nbSJQPQ35bnXSxdqMVjVtA05G7pnTZZOF4BXYaaGjqP/vG39sXTUtwnNl
3ZtaHRM0tYQLqDEXcErAyb9NhgFTrZSN+frZS8mRNAGd9zTNR5kIcfXwQiHrQBEuA+bRQrhOGSeX
hOSajVlBeeZ44gsmA7X4MGBaPGxBiSbcw/EHkFt8qI/pIPyjPZZQUUEuHv8N2jbY0MTnIXZ/ScrL
HOSuBVUOFsBkY6HJFSxB5ZTXz7AgUAdTzuRcCH09CEs6E4uzlf15IXBYe09vsFrKZL4QmSX5rPbc
9UyBprsHvJjRWvBLX+3ZwjrbP5kNUwf+Mo/H2lMR7g9wxPEqqQR/w7qZT6Hgk+kACm3I9aDBHIvQ
FAc0L5kapy9rC45PEv2UgPFzopVDBsU5QzdC4OeEyc44IBL4PS451VGAp7uei0G2pg8eA1L/0YCW
dSfrCDaIjeks+j4Vje2AJs7fJncidLetIpc01yf9VkD1BkwFQwdejnpXFV+FzQF9/Hd6rXsiBrd1
+re6k9GU6jnHplPPlMlPbaGyS9rlhJgg4mTXZjncePjLvPAFyt7fn2oVkT2o9X7eIm56exfHOfKS
56Smvj5o3jFmWEoDbjjU2RN+bHQyfk0s5uVYrEpjow0AXTkZoaN6s+rK5kZWeq/GBDJWV4cjFd4Y
nTpDeQuQbO3B1ttEOCbEP3aAwdrg8GoQI6G6JWoViRsJ1GfWLpg/wyAfzFg/A0XJEmjKzolirG5h
65IKp7OyFUqgQhY0+fChA+mgVA5jXQCxBJTMB851wwUbJ4NxPtdSA4aXNVS89YeBFtXqRxWM9FSN
20Ayzca1ai7VWuQAxWbbNzxGxNMZJWWBS07BTjEjD4p476IAQYCKbyPYVq/WlyqAmdfMUi0GDvaa
3xrj6VQ7D8fciQBiduSBETVEOnNDx3gGvdscIdFYS62s+cSGjJkpdRazlsPDG7LKqWUTNNkwyUy1
uzJ/gM2OBMOenPKHNT3Knnc4xqDCCK7z9kkmRUWmHsvIYYrcQF31BoN8eOG66UU1rWunuLN2fxGN
A2b5vzROjHVrIzRDqSTJ1B4HqFDvLi6IDrf79EfcY3DLnKHCEqgnI5MsyhOMDPA/4lSLkAqzRUWH
6QD5s6TSON6EYH/pHkutjGtMNKfBtiGl+wyTcIlwucpBX9yd6yES8xNJo2Z1fHkuEvvkV10zIboC
H8E9wcAgDk+75WY0vmmhOKXoy4JbpNftQYNGYAKOs8ynruYDgtHI6qpcL4G36q9Og96CVKCpVFye
EW1xCFb6HSCdDwO23C/9rra8pnzoQXOzuQ8Gc4G0pASK3tsXW/Ldcpmu0KQfbDwsCJj3GZIQsA+J
grxjpfz0wIxe7ixh4L41BF8ynY6rOdhHZQT2z3g8o9n05iBl457qCJ1UOA8656T/wzmQcIm+q72Z
MYIUGJNUmMhOw69uja4487KGbn6NnCiJRG9AdDRSx4WaEuoHvtvWW4c83W/NgbSLny35WLeRDzT6
FvP4MUFYyVU44+0UYRSLoJtkdJ18egwzSfJybf/PdhoXNbCXVYQkDy+tM+Ai+sTGRUc1QIGbclgM
OeMoQXtyu+leNzAWDsY2FDc5a9rJnHYO8cTxDvCrizRJqBcAVn/JLh41/2hqbnfN2k2dsHpW/f+N
WrBYFXFrYsP6haxugdFc8IYoj5FL/C7xPrlSCbc1hYtHIf7XNE64nk7Zc9EG/6r0SfRrI7M61H4l
zbwPjLG7qk7MuZGxVcOVf9az8n4JSeTezrWFqhI2QpQ7dm3Jd+sUgtZXQ2bmyDy+EeH695I9Xz4q
7KwZnFL59bCUcLEeVl7FnpVs97ne6iq93ZqH4kvu80mWtNR69WGmB2Mzp3BGnsurXbBSs9DP08e3
YwH05zKBWpgG8sZTU0DTF81cVl+A7kF4dU6Fco47ehdhI74XjsMA/RfKRPlekGfeuQoAfbtXScII
0XSFjZxpzE6pfdSKc9bCML5MPrsIppbxMC1sotsEGbjh5z0G6ZMyNqKlOszCKGIRiZesMf8gRBVz
46fzesYmMpcZnKNl/ux+pmDbdM+Hyx65WuUpBb5XK6EQ/4/3shTJDZ+/3XFaTsqzrfw4hnDn9EMM
tQUB0n7KTA+lgDWsnasFvEgJq1PyWCC01j/C0oNVXEKyNXR1XkiKl/y/HUsMmGB1RanCg9vjyMRi
vMCUAWZn5lF4kZ4KYQsL3DivdIehEh3ESpCQ88K0H8Rs22wZxxIWFRdHwO68lpAniSMZStuLEmcS
Cg1hTG0X85gPHWhimb+onRSI48r3PvXYi67jebBFTPeblFzvuTdDZCp4K0zjUnCw0HiiMD78OnK9
aDWnka+Xo+KO72l1hWOI8ZdPtHW2qFED0dL23rHouRyVC8/WDpAZvSaEsyk0LigmzW8EYQQjQTVj
5QPAZmcGcP4DnQOpDz3NbaaDAqD6FupMJG3XLiAeMu/O6XZxMyoKQjtkvWneoi5EFIHvKejt1+E8
VneyfIBVaUrPiIn1qfHdF8h0OfJzkm/0jjmuGTct+o4znLREtVTTQGF7T8QJwLxwfe9t8p47E18E
YG/OJxrHpndumBQ9XEX8YRbeL76KOP6tICE8VlgTd2Hmo/WazHiWyiHAChSnyh0ze0DQG9UXAE3y
Xs3Jzl6YGsQ4raZ99mBcF2+nDlMpvN9kvuH75lSQu2D0VVx5rbJ9Ekhttm93m97e2QXoK2OdnJOj
Xxe+K6oHu8fOsfkAc17Pv5c8oo+ZSsRyxWpr+k20ZASzuIEzqdtgk/i/EvqGlkihWw4suRTxO0S6
B0MXIrWvJrAvHPL+7RYEs8X5McwZgq/MxLRobHBwHCpMMtrht0slYSRaMdJcTGTosgQ7FMaS6AN6
BotVMHJedfQ7v5pFJve5rSepWm0HZwcmZlKrp7J6S9UesgKpGE1Cb1klu9QlLbV6QUI4/JuRqZGg
8BNsM+ij4HkBxPcBD7+Ez0m6xwVUI5XEbeoxcZ8B+I7pixC9YgbXX9uvLk4XNWqauPZjB3FNU42Q
hsmnddOTJr2OA8EL6YIXeM3ZTpBSxx/wPr26r4pxE8V+SRWM9RJ9S3fE4rGeJ2s+jUIhdvecmyi1
VWecvo9XGcMIwhyXJF+3GrKGXzYwm2TdLT0bB0wFXJor0fRdFzMG5aGeEmYPUET/0y5TZ2hknQ08
gx/xCCIIzivYruBSAkf1jcjnoF4x7PCFX2DqKLAc3cxYkIJe77yaLze3MQ0Fml7PH+WK3Buvo4/8
ZlvxQaJdMobNbhuB2XClrKbtnxgkC5NDREl6xQFrG/CwJ5H+jhzNXJzUBldWJ9Gb41azQowLUQqG
Y56ABjjam/VhnYKjIPCUwTkm9Jqljp4+mrpeKxHvB+nts2KTyxyk0xNZyI9Ls9R5iCsx47reyZXH
BEuO/T3Q7Hrxby1FPgumLF1HwJxHVLFJV11cBTWI+53u33xIGeS3HtriGTokefbxirntzuMPSaRd
EXz0MGK+6WLBgDipp8BWUrdQW076h7TrJYIuvqFX/WSK4ljn2jXt/MsQpGHEMTPB/st1la0BRI2n
m+OcEoNi4tQ4yTi5oWguVHDtzXzPF+l2YjacSv1p9/36sJYVKWUPtvNNM1ic8DEKTQonEGbzEgCY
+YaEdlzl8qvkRmUovpnZN8hTE9UgaV94XTj2codxkr7TCW9f/VceVg6oTBqygfH8YLcIXsSrkxeD
2ZMumOl3UwwcHZAJTWyesVbp/1UbQ8ONA0OWz5FDX5aN3M9C6GfZU+sPFXmXHyxzUX9j1zNlhEY7
dMZ1exagigWg731wNCg7mFYlO6DAo+vA8e+3n1lod/tcs9YipW2dymK7vvV5Q/K2mWaSGDY2MRP8
zlLkatiroasmJVVdMbILl5F3z39vHT3eiatvEikqOV4Nt529uENm7HUisnW80XqoWNZBc/4bc5VM
CF0FjJYYHaYx4nA8aO3hQMvepZHl6MKwVk5jP5kqYWqsBcYwnShkJh9QPKIK1lejNdIOhaOSdST+
PUHiI9UGcNmg/vIu2RK1+CDEtlb6rodO2Vq6g6fb8b2ALVnPICXOkL6jQmFIgiyOpXGbPYZBiADr
J3/09LiNjzJk+vWGs41mqLsLWHkvFskyV3K7VzC3w/hPqMDLBcXnM9HRs4y696a5gS2vlv1eJmNr
W822j2JJKzMVQJ9ky7Y0n6UJwlRni85JKOh5/E/hDpkn2Qq9M9bIAsPEppNU0dhAmCUZeW9fAj0r
4MotMigJDzgXOvyyTlfPt8ZDqC66iiFL2jRWzHD/aG4T8e1hpBvOqOMrZVlN4o03zYHVmALBNY7n
rXpuokMeiIdAMOgm6H9qqQr4taKDze0EhnwDYTCB2L0llnY2Se6TEXt5TcCZ7QI6EyNYu1Syz/ih
SsT1mecZTNPJDEdEpLOGI5rPwS6+zZz4/st511NhJ0LyEpkI14mw77maa+KpcPu303c4F/vWyIP/
Lda7bM4IgwMlGYygJJoK9d7ZoU/J7HzP0VKAKcmhUyO4vNIE3M7nqTWYgbbyPlcrUvlOGtVne5dB
x+31k02FQ1N3lOx1ZRhkhbmElbfozgscRGjCLS67s89Um6II+3uCcnWOcgQLpS6zvT5Fmtk4fLca
l0BHzPKDY2/ZlJo54/oOsCeIwPeYW5KlqD5GlLUoqIbAKTjkzCzBNsOuX/XRRP3aJvgENSccv0Fc
+jrD1PeljddOuZRg8SVeX4G6hhRDuh/v50EO8vmC2moy9OnY0KONZeBGgOVzaOsJlmsxPKA2iDVJ
T+V+e3aictJzcEcVXeibdHKs60u7dcT48X66OsyRfAdm0AOiA3UPWRrZE0N5kx4DLtAw6vqOfodr
Lubv7uzqhaTULST2Wb7b3NV7ZcCG1IZIyWYRI7KAG/6FvQgFzD2nPJWxs/gazNF6+BIBmZaraMoF
6fJPX1DUnHkCuj4xjvfMf17q3tCWU3g7trylMIDtiUI4eF1EdNbI9jCtaLm2BAf/vsWxq/I8iVNd
oDEdtlSdxYx4dn09oqLh0Phylv1qcHyXzMt4J7HHyC7Fmk6M2Zf+ilyWIyHSKVggJoweCXz5UISG
8Z7sJgnbkdK3SiCv1b3eqUeyrNOTVlOWGrrNFUEUwTPVyx24Io9VsWpnEiHN8nNi9I/HoVG9oph8
MlIZe8h8MDGSKv66AhjA6ffrmLRrbNypaDCsXl0V68/Z4fTfqrmQsdFEYDhJ9f33zGzGjsIhGwG6
pjpAIN20mmNw70X1/5oIP91mzHXnIsASPgvriqJ598QbZy8Myfp4s6YEJji7aYdf6IA5hvpIUvfx
ONwpUy5ZgaLb7xbezb8D7fQj3Zoli0yWsTdlSXh0AWgtiT2SM+n7DJMFKDbi31Ja6gXRQL4aSYPp
AdMs2gUGObNNTobYkZrjvcqJT6W+/EJSV4Pd9iO7fq6pZ/6WMX6LmBLQGlzxg3iRlC8iGKE5/8cK
8AXM5y65rtRvP51E1NOX0fto2MjO/u8YdW5DWBXuyB8Y6Sgx6ubFvfOMEv7Hx4frVOiweTX/L5lZ
5EtwQwR/W6/jlVkR9h0NWTiKAPr7hGwamEImnN/d8//hhcA7HOI5uAJDHZcwwJHanyaT3rj1Z45n
+pxNwL6t4hRppKEWBl6a0P3sR+PvDSjAyN/xP672FMg1dXs65lxYeRFnSP485St+aOjNlh8DSK8e
2tfto5N7ppQ4zQfdjTcsEE8KMTvw/TAEBSJuaaIelqyGEL1IsPEuQ+kw3Kcw9GGCDEPb46eif7X9
Bp0LifxRFPExM8Stg72K1SzA5dsENxv0P+e/I6b4oZ5MkkAoesJemxZBZw1JdaKYfC/oY3HLu2A4
CUTyfyWVopcCDK48Ye1xZ7Oiu4sWaPjPdcYP+4SRYDu0XsFkDWaRMoov6DFqj4pxWgln6xnvonTU
+uxpY/FtUsMV4oN6b13xltf7vQ+Z9k9QGAI9Uw+g7U2nU1qeZ3kGrvD4TwSHwSAAYWecSAsOk470
Oqni7rntJ0G0bTtk/70l5IK0CxH8Fe68YyqbkLQSBsaiZ0hsnBVpOdiuFPyBFZMWOFb4Y7/RYQoO
DMR9P0UuejrcInsRqY60f6PJMrSQ295SejokApxpY06rWZex6eHBgyS3gcaLyezzgO5VR5X5wNTq
Pygxhx0Ibo3aIaa4hnrXVXFgY3kc8MrNA9xCvdX7D5qEmtOiWh/Fhsr6dvjysrhhxidAjSq+37ME
cJvqRxrEe+PjM7NUX7NZsOXPChmXJurCEG2KgDc99FDh1FEjXf3zoqDq+1+zYxA/Ol9Y1vKL0946
jPISNvLx1YZVJHEJK0LaY1+kvupotBXXL90j9CE1B9nkn8ngFO7wKdPhhaioNzS5HAAob8og30YO
oy6/dBZd83kzNoc+4UBERruZWVuWKPUravI1sjAr0f927PiI56rc/nLNBIHuxz1sBhdmohmgh0pY
IqtBQlXeAYX3Mic/z+1XfI5zDKZKTLGtXhSCEXA8O6yofRJoI15DDFEDm9WxH6hy3zh1H6cy9pXz
sQ7pNeaw7DoSq7N+vdlfUTsA5QzmTJSsh1BHkeXiUVOWhRZVIZbvha97nxtzEAUkREfhoeLE3Dym
FX4fgKVFjC9AwDMntQc988ssen6pMYttP8QRAEWEcLCLmd/kaCA3Dg+kzCSz03xWEJGeSrG4wuOf
6lUlJPWadSFLsJH5kjUqpMnf25f85q8g3vXJVFG7KhXSvlf1t32D5MKCQ4lV2pkWh3rFZ/EGFv/d
jAjNhnhuxEkp/KWx7icPaLcH0vloQ/Zu9hm/pA3PEk1ZLZ/LBV3HGR4NusAgJKnn3Syru+qE8u7x
25cyUBNaKhva6BcLmNk+Q3rxQCFZYhfvg0J5+dvK1z5mp/xc7z1nKP9pfJbwe4Z3sVJVAkyGxrun
1edHwIJcRvBYcxQlwl7iE12pLnq6mwd2zOs1RdvwxKTsLC6UcmPtIBYNPL9UV9TAKgFI6ezaPE1H
z2bVu2XaOcV/Owz4zNyf1P0lBqyJb0qFG7hM1I25Z9fnk8hLePIinZ6rH/aPsLG0psItBhUYXDbR
To2da/3kqlEgqcKHsZsjAgHl2RRbQsdkdGpmUbmXLeGeVRA7bm441sKDubAypAZF/oouvgWbnQ/V
O5AG/pqWvo9CYrdQQyPFiFeYCaioipOri0Ey7JMIadV13gVYzL7bmBawzCy8lClv0U6JnjDsYJX+
sfmwlLHKMrIgLd/MDWwRwMyDIEWxT/iBRJhyQbAyoqLfvN/Xw5GWxqlIITejs8j/8PCR4aLSRGnW
pj0OH637cN91A/5IWRVu6IEoUhm0CNSS6Iy4PQx/z6Xy3Lqxx5IYBa9UaViPyAJr8EiSjXa46CYk
q2+Ij606oWCUfBOm7cFkmf8HW5IyKuOY1LO4E2PwE+WS7vyclLk3E8TjjjjH0LSG/Bf9+2u//8SR
UY1Nk5lne5U3ETvGw0T99iMGmPRFfCLoh1SAQwBL3vMc6e9K/KK9L9tCRfoiTmgbQaFIJBH4HnTD
rCxX58zGXF+5TqskGZVqdkK+wz11u4Mz7LA3AkWzHfy7sHnbQv0+fV/qpS2cuUSjlAoy8sMwtafu
DiF9eWRF17ELeciDCkCLgZK7ttUcjFFEJzDMMvrqpyhDzdE/I+vjqeztgAa4dcKQaAGMIWvm2wVj
06LEaV5tKEKWe1U6OmVnbCe+RdWuUjiVnuTUnBlE5OidywGz+OJj6xtdEIUBJ/BGnEUfaM3ME9OZ
sGMaOWmQwJFDweqEZibqU26yx9hFu+TpmQ7IFA9KQce+jhsOOX/OCXesBOyEBIA/He7NIrsG851y
AtC8jla31J0YS389IfAEoD6B98WVqTZIi3s/t6bh1MAGyVtrCxEjse+54sdEA4xRUUnb+/iyKWRd
DZtVJQEUt3vXXTFVW+N7ocRspqHqhLuo8PoWRMR38enyy2eUaAhAHxmtoWepobARBA+BnDaTwTsy
jYsVJaM73NlmI62VyE+SQh/S0bDU9K3eH9eddBFYX2KRqY+/YFRhTtPqmipK/dpYl52DR4wj/j6l
TXEndGqXexcJJ3xtFvYxpQt+n+3WDaCkISneWw/mt3sVKkNPccVHdvi1Tu6IkA0bY3NG9A6lz91l
7irmkTjUTRyNnLrzokn1x9VcypSVe0hPDj9tfgVuqj7FvvkyntHMNFDJRH0OR4GcSyuYQX05kEXa
kPTj5fi7GhIdOnoDRa6XMVf1SWNK1VgWbOS0r3cSB6LhR+PewtaUZu3y0KjwKKckZ5uL7E60aa79
4X0CnIevkDlWV/1Fekb3qmCMSJA5HTWCYUP+RbDAtVMFDw7XMzYDKF7CzvtVJygATKluMuAOQzv9
lmstO1iwrku2wEfacrTUEX4Jm5LefPCKE9fEtvYo4OGclh8UxKN8gGiJP4X4dBXEVq4vAeGYLEUi
5oEU2T4cn1FC/0ieQBoab+PeVuMUqEOVpw9HQKGEEJf0aCg/AHh9jfC1nOi6IMLzm+OWYtJSXd8L
fOeX0ggEfmG7BYwfTKS55W3sQqTzgkI2a8T3VWoBKB4i5emoIDUuIYR2l6nr9scHyp2oaP3CEYQQ
Iz/Kly2Z+wVdRnJdV3dvKITr5lC3QEeeLcmBmSIFplFURT1PHB3UrNhnwgyURPvhq05l7z55zPPL
g6G/RxrRcC8UbdaoKSPjIvdMbf69XJ6oqZLNcbWrM56CSgq2ajlakyCxrSaUhDruCFpPEeu6RoKm
G+qmo4yBpX30MOXzY9XeMKPUB9WJYisl6qZPE3DiRyjJo8clJJlU9PD6epFQCA3zqIqhJWm3Ub/W
0DEV/RBkcWi5hOhRaIeCS3Q2a6mqvMPVopnxDk7oR+9tML+sgSnuCWZt5qJ/JGH2XXOORfvkwMVh
SoZmbCn4luRVui//3V+fNQg1pj24ozX4q35UW+p+dbZvsxle6U2sH7wKviu+YbgL7t0w/qTcskra
gNJhfssIpweb/g+i6fcHjKeHKd+LZHCgS5ULEC3NfPi36YAAhSAy3Hvp+1qHKJLJZnKDSmMnjA66
V3eEQP1coOwnMkY2icXoJd20wsdgZrlez2bC908NiQ1ufDaUN7muHH37uwsAU1DLZ4c9L53HZxBX
9fzCFZzhbLPNm3m74Vp5RQftLJl+8ixB7cA6OjjWCP18gOTJPobxTgiDkwrUCpqf4HQRq3n1vTGn
LNoSb0FChuwJYIpBvPp1V8YZ/xJrh0Dp/iv4pJFm1DgsLTlYd+ClUlCYrYrNAWYb0feGmYyKpLKg
vo2L2olJ75qW3UwvGpeNqlmPHJyA6M9Xl7wsUxSg3rvW2ydxXYsilgS5waivlgweSthtpKsPn5SQ
XhivJJ5+YKtLK5GhE/KujRDkt63Wl6U4rV200VykdztTdCMqt+s0jGtJ9y5KY56bxLG+qkvwAJT9
LQOuwbBC+qvXa1AGaYhEzsX8mGJRLebi+N/V4vLJkOg8EJS/rsacFUdHYN8zeOdO4VD8RptH39RY
3gTVXb2DmOJsVGazpONjpdbAzwEDf5CO2bKPII5UhL06vrrMh4NhzpmnX/N2H+S1Ke4xAGNdk1VE
s+AqK+4degrivwxV8yOsUT22EPtFF15tygwapZaYeYVFW34SC4ScTrLf16ZyN6xKMZNcaAe5Z9Lm
V5/ls0WlvzsMHNw3szrSuSeqRcBpAAI5qRTe27tFP5oGC9nnT35z54sIc9Wn0tqWJgBISiRb2plX
AsXTGK38k4Lo0wiD28PZxD00SqZPY0AqnNjzFyCsedSf30bjs/yJWTnZtVqktsxcBOisNCvj10mL
HCnCfTmPGqC3vjTRI8fw50XqHLcjemlCEYujiKw7DqPtoqmEmGpMH4rNsARB4M1MYDkQJQfVgQmJ
XHhqHIAat+6ub1ttqYS8NPXKiXyrUf1tX3kcVERfrporX/vHjyTz8PS+utPgn1vq/AWZmi0an0Ib
fsr6maR++BmhaS0SIBIp3AnlgWOBRdnMdFw2zgz2H2D505ywF/Hto6nvBKqNP2CrUwGPkrg2Ri6c
gsAJbqXPdLFqXzkTHItVaboyymrDvUDO1wKcz5SuoqEpVXu1m3QAM/ZX9KDzsGE6UPSEA1m0Ysz8
rrIMyzcCj1Zs7mTVEB+LcXHoAbK8IoNh23kg8od4QjrDHXdsRESXUHu5rZJ7V+syR0zCWS/B5ely
wZBsEMELeo+IAMhrhr7lMlvEEosjY/PGwi+VsYeNaQv019Q9QFQG3rkQ20q+HPAnzx3W8YHXZR/h
ZqrWNSg9+AgWoitF7c886vtJM0WaP2F9IduQnEMz5GyvlJpPvXLmOGZVX60TWgiATXGnbPlJ6F3l
o8QCeXe5orWRf4vCB65iyh0dUg2kjiS8ydWr59p3iEiyp18Jl82uZQ1Oi6K482VA7UgtCqnireWl
iHDcT4MovJGre7Hi4W0qaC0UOgghnVJXrX7kRhfesghz4gyvuaA0oLxRHWSFuuCZns/Qca3HPeWJ
Hr8qU2GLIDkElUsdrDUVRdy1n+6MRsXBnWkiaiua2oe5mMhMNLOy9lAjc/z+soJE01srR6qBrpE4
6qrpgVczeK1VYaG0+qs0fiEplEOvo469lPrG4odUrwrw4wp5cnPQPFS+rfbSZ+RigAu7Z72yi5Mq
+qWp32KYSBw8gM7vAcuFyOR9enqJLLqO2mWHJQ2bMvVYsbRAN5AMPXrCubNxc+sM639Oi8/Z2MuR
ygDD9KJ/MtZAiLZL95L9M9Xt6K5MXW6ZVjg6X+Pw+Mzzm/Rm6UqzpskNtEiBK8gbE5iuiwH7bshG
MwVlcKTZOV4JkKE4csf2K+CCtpeF4yl/x9rhlGJNKltaNVRADft2gYPcakAuFGiEOCSBeVlyfAoq
QnxPpc2dApFC8Fd1LPwMVGEPAa7dH9G01wcrJsgiv/BKoG6er0fcVj3pAI4mAW00Inchq51k45Ya
kgrqemHWHHsJm35hvVisxeB1mdOuvTeDtGAbkr1sunBgExDTrPy9UBykuYR3J9GelUDcAKikwchN
KkS0x15BPMEui6mE8dNh82+2vmkZj28RhdfiqPbNCmFv1n+tE1Uz5UmXnMGjMIJzJyXGaj8G5jc6
+31pFJl6TMZAr5KO9JTxO2nxBinjjkQzVQTloXcQn+MYDKfDjLGlff4qK/MZ1kFsFU2vTvwJNucB
mqqDW5pTUTkvhQapsqSxbsIruS9JV4XXWxzwco75JI3Surb4F4cJuLz6PB9e+7hcu5rERNoMhbcr
yt/84OMVbswoHALl3/KM6PmE3qpgF+ZDG99urnpjw7JJCobIFrTh0t1uebo0Yqt31kDJx/0Q7rDJ
gfCgv8/vQoTpQPOWvxZmrX74LIplCed7KuAA8T6iz9JYavctk0FkSePz/0IuUXT7+koE52AWBK+T
I8vFvO2VNwgOavO+itayBqBoXsTNRbYgRNFHflL4Tz7A/oWBF5wUzHYfeDpY0DbN/XjUEzv0CvaE
ub9OYQno67q9FLwBhQ9XdMEIduqrmpm/YRg+jkFRsq4o3+Vp/qyeJEw+vi4nt05VnTqiSlGBikF9
TU9vVpVuI5Ztrzal1AuZ83XGhSsykzkMKhGbcCchZC8wE5Szauq+Kvm5kBQ0tmzXcIpjEiLUJwmo
YY5ifj8CnkMLxQyVN/esq7K+alwXnKRJxRp3doM1JnADGV5n7ki2z8wih2CuLiTvALO3b/knlO3d
0SZCBZXR1sUEB5MQRJu0xSjiXINjkxUpr9nHcfHLo3Gl3NEoNwO4eYVTMVknjg7I+wgSfUQzNt++
sQgSZlaB0faWCJ406LS6jrFp2d1jXdUd2SKA1t2mWONRyZodsUpjR0k7cyh816yA8b3bFs/9kKuc
lCGcaHfNgDiV3NDT+rg3rm81i2v4nXmavkwRBbb7bdm4WNMLj2h3f/kdpWUGJYphQ/EZgkO9uEgu
AWKxi752AumVaBr7l5RIIzmDYbRv+hTipF2vI29rvZGgaEHRZJf7z62HG01qBfKA06zqTyJBglKX
ilEqgZUQCqne4ONZiBeWvLVKpNARlJ2Z0auZfZmw69yAWcyhAjSD+nBc+8hCjjdc0HDUjQa/eq3d
7jINBtZwuDIhvkZv46QOzP4CD/PXREqHCSZRVQZf+xTgUaBObxc5rbgVUpViFNQiLn1Lf8AyptwH
CwSYi6OnWOrczvG0VXLZ5HOfaj2C/lwW3vej6EGZPpt1rbL0gYBBpSchKBOYN7dT6REK3QLHvqnF
hdsUVfGwIIADx1iDuqVPxyRXPaHxMUpRdgRFTvD4D/RMrix0Tq7ekIBgUen2ZjuOtWHIeXjpJ01w
xsoBqDzKJwIq9Sw/5EnpE8FI+T9tKRsy9NW5/mGJrQN7UCR+xjXxmDw1/4AT6o9kD0aB+Eh020YL
WScS17aaqIOUjhXL0CaillDM72+jey3O6mUzHLILOyXyRHzuTmeMgihbJnWR39p9RUsDpPNjvC8n
Tdcy1kUxCD1PI+mDiu4MoYQqW0ecsjlz4Ujc5msKpVaDFVFCsREIiwI3lJk8xMRXFC9H99aCClGN
tNhKk1/wGPu4MmKRIzlHepqEhk3t9VFp617V5C6HcMYTaTxB2kl+fLX2MAZ7eM/LaIwhdTt1nhyn
Rq7XQjumOuNkk8+9G7i3ct8jKVCWNbtW/yfZ/OnIdAMLBKFWJlbmAdR3symATONbmHSZ8/EQGsxs
xKK3ShBXK8K1Nx9w1SzdTxorwP+1WYZ6KW4egIbd90BPkVl6hQ/kkPJ6XM0sUwxVpllmmr+Uq03t
ABFEF/vtXAVzbuzWSHI8CXzxXlNSs2fCwn8rCgz/9waFmz57/wRMNGk8aW7OfE+gN/UQC9YD8UWA
ITL9CSIJNK1jmt+PwmSOPDXOmH29buga8YDbwIpuEwTqfO6685AsJTBsd8HavMAAmRhDZ/myHKF1
dyLImO112uM19vcn3arNS1yK5rx9MBq9qsWJtwQwX/lYwi3PGuxT9EWXw5orgwwxM5/7iE1vur7i
SGJKiaPyfI77V7rQ1ZIj9BlPZ12u7FZk53CJVE7DYpsEEFFYvuU9yNc+H9PPM3rCkgSB3G1v55Mq
g9mLnih0c5U1rKgFPSIJGCD+4cDiIjFjDdHQLdZKEetOu/wJCuASdZj4Xt6xS2ZYfcmjzHveKBu2
eSB++rhN5oDTNCBbF4Gj9+zuQ2oUDmcCYItCAdr6gi5LueXiOVGuNrwuO5cRp8oEprkC4GzU5tjR
/zCYyBW4N2iIbqQCGwVHvAtLpEJ9Wiy98+Bq78tkeSBbdqicjgbAC7nEMzsq1zFBd3Kdq+dXpmUx
dDZpoTCwuCOYb9Bui6ku9NRq2/wweLEUUrSfC5HWNoqVpFcJf3eThSjvJI5XMQnMzgFUcgk7NdsX
vZvc1DcNAH7iC3q50jcujfgSay4qPzp7PlIyvZpxbbiubj8mffBW8aHK5aeP4EvF7KdcAhinHeNV
NheA6eh4HIQenJyk/PvT8ngvuWPR7KuOyCrCrQnY5Eps0Xh5BQHUHiCufE/FFeVc8lQEVoBwoYVA
7ulz+y/hasqXr0D6u0kFGVvAbHjjKhA5gpzNDaZCjpqjuWI35TMJcB4GMaaqOUXKWWxFI+vgSikv
Xqnb36RI/YKgPd4exg7Auu/6YYAoGWW5VHO4nrTGaCJtkiP00Jjy+93MMtuVDe7TQ315O1NfXEB+
EtWB7cdxc9JJu6/uV0oM8Qg8AqR3GrFzgM+fk5j/Iw7zQj+hm0cIxq27FrWvmTPNwhNlBQZYKxdu
1q5/cGXW9ROOYZqpshZyZOcEg3x+G1BY2tgFZRts32FKYlFNmyeyAKDU4m6hCvIQ/2VhLdi7IIA9
5yUq3AJKFtRCzlJA/d2QfaAJ/3XUPuadfbQ9Uz1vd1gG99n5+vE3bgaPpKtPfclkY4Qr/CR72AuZ
f7wpYhYRotvcaFcDyBUmwmi8fbFvpnoh5kogFtuSB7NFQS5yGTbJahenh5SLclmWdj0KYcwHSb/j
JWpwr98CLGK84Rl2oQLdUcDOkM5Dvm+AQxxm9cX15AXGqV5cErClF6yp8GXdCf68f154JupaXQk+
yvwkQdONbsMKDQolb1k2jIGzGmKbIWHopV2kgqAX0X5EoLHCVl9wrHqo9kRk2h5mHO9tEoNtmuMN
TY/hF4VVxxrd/vIen9SBsooGEvguXYpPzWkRCEQXSeVtak1io/NAXltnRj3S7m4JHNr2DpDx9W8V
2J8X4VbFLVhu0NsSau42LDjfNlis0l9vK0EvsmYpKBO0Wr1qWJWWG5tXMlxLbCazPIrnY+5J/68k
cvYaRq1bqcsNPrV8ITn6W5kfP8atL32XCi1l+TQwK3lZnESKm2QGPHvBl/rNcFCakeqRTUCoUqsJ
PiUZ2R4tHeU/iwyzmUfM1OIp6gbyEW8zWxs4L2BMl+mfjo4Q2F8nBWYCXUhee2ORBgrjsug858u0
p8kU/JScDGh16oVVjtYlq+ZfPw3SrMJG6mdLHxcqtFulr79kuyfIpFdCbirnY1qxwcw6Fh2+hpKa
F7fh63nZWCzNLnC2Vl8Qna35YxGNoH4yxj5ssmRohmiu29lPNxOfTC/EoIuGJP0GiGS93Viq9ZfY
ifILzhv7D4F+VuaEZtluDKBzXCI6TwKw1nZvVU5Q1WkMpSZ1ez7zCRpXeLeniRDiGlsMXlXAg6sb
Q50WNrLOKx6btpBrzh9txEX4gIMmX9C81H9MPeQKIb3udURDqVKTBPXEYiFFg33RkW6kmR7BcLsb
OFvbaxVMwnzRp2wVF2HlpcptzUDH4RDjeQpq1eG9VuyW3LBCkTehhOXTYLK7LuWBlHvSO7UC998I
nzjvHfIHzh72DLpLOHD9WrJn/r90B65Z6ETDXrPx8JyBBGMgMntAewDFIsS7zT5Tk8iUOUyewo1N
xGBVk/zIF13aMFxTj5CSocIvrpWWFRqb2y919mKaM4Vs5auon1dsbCThVG5ChyzCtBETiDy1+8an
QjYczc2rv6A/YIJd8vENhTZZZCjMa37ovzyMSkhQhXH+QaFHzKMogWeqxyH/gOtC4y5IWh52UB8B
pS+gXMKcjb9u7bsHikk2t7Bfl7AKO6XuGO9reyUHR5mo5d+60l8WX0yVgf29eUus2Zxs6DiUotmz
QmGefMD3YaJLn0s0sFUIn2PRMz4mdrO1iL2cQhqO5Xt4th4/ur34Rxc8aAHorbWkKLsibImWbwgY
VcMrObb3QcFLSY+938l5CvTEqCzXmVq8fLLodV69S65as+KNVz0wYWU1I8QZW2pGwaOji0QkCfr/
xT/2ept7zB7h6h2j3qtWGgrbsYOeie4wF+3DrSTZEeQqKy0Cw8qWriOujv+9FZQfevk55SD4H980
X9+mL09aVZ6871jC7U8puE7GEekHSHBMAHpecXSMq4G/UaSkrL3mqc8NGVCYx4BJA/6rF1rM2/3c
gpvQLyN7AjMa9JtU+UddzhajZUYnOUk66wV8XB39T429EyVF83cpdD7mqdRgZtYqrht+nrPALYjS
hAk8DEFYNnHzejvLreo9KQdNyV240Qm/FPfMFTsL6e8iLSf8AEHasXa6fleAyh8y1h1JhbVPaszo
fCohDe9c0LCrOv3+CO1FQAzeABcnNQKZXa+uZhTjdmJXTD10s3O/grnv9W5wbbcBM9QjLYJgAjA5
nP7N02IHTMx6ljN73aWLI7uxNeCs4TXk5qFtrLFeYazOYL1DTwFPBI6O+sz3g5T7ZGYg9Hwpf1Fj
lwYuUJYAqMq7h72lXWsE5LAF5bPxK9l95Y3c4aAW8a7YWccvJWGUscn4TF9x8cvv9XnGFXLepB3A
uPqnP7IU/Gj1fP2O+X9R3kEJxGFwYkBqCXMkTA7y/+9KIWiowu0y6fezJclFfoTH4WlkRwtSGZyS
n8J1oq3eOlCH00d13t015vwIZK5cMAl5mDxTykl8D8AsfW6lXZ3aYOcEHaH9XQU8Y5u8C+sGmUxb
MDrllYx1JiMZCe5moF70IO7l3zYw8gW5/7MaS0p2h/PT1brniqgGL08OsclK5CjH0/rTqUIcS2BE
dHLsGeGXSDy/uKZsiVHjwpk9P1RcL/5sMndBCQp/nuvq+3/yiW6z0Lmml0eu8Z3jVvXmIPFAAhhD
+EVZ/Sn8L1w6qtG8/7lR6OjCGzru2G4yItRNaKbIW1seYrKY2rt/4mSuLOPHLYuZyInorq16XEDV
ljUDoiYiod3l92vG5aWWMraVraLMR+++XnvPfueKprdrYNMYPuVJIbePmOADh0BgbWACTKEAJ4fR
39on9ZnWsDz/HE1ovl7mywYKxCfaomK5cPLn0US80mXdUvUOkcqhjjiCFKBHpyX/g3U3FzXkCM6J
AKCseSnDOLDnWsLLoffzH4oHT74yqXJrRld2nD+/brfx5COZqZ8BCbcK+/4h9BN3gnClSV1r0L5u
ZY3tVIx1rP3sAl7g86ZmTPlaMJQ3btQPbIL5YwaxDAwW8bN4wWQbw5avU83YWaN4snQ1QBzfKnZL
sQxTvQlE+iskaavv7GpcyBHKKEXFvG7aKd1NFeulK3ZbPEW4zKf0w86aj5PplXOjDDMsLK2S1UlX
F3XqvwmU08dPEc1vk0RLjWan0hi9VaeFUJ7oKYaabzoosOmJBGFZd1/IIkD/HlQUUlukNI8NxSYL
cTe6+nnprYiA+18DE+S3rC9sB8WUHgzD7RSZsRVrrY5Rb6TSc4FlunOvBT3PmWbW/Wp0lIu3PsDs
2dFhs6Cq8RR/gk/npjMlmtJGHsxSXTuCH78LF+PBHXJ0WPi/rQM1sknJu41RL51dqZr20BgmXSqI
W0u8SBB6sGIy95apvM63ew/WYa35EUvhSDEYawEFrGCP919g3bCcd4jsVGjA2l5BrgQRAC/5RQwD
BeS2UIdLwIiA3OYJaOD6DYvvJDwQirz3m25FGjnKXXfinWnTrg2daYV+V+at2fm+czoyBqpTKda6
QdDk5qlAjBgJemSezVy/a5XNvBoqDsbCa4ZC9rXfGkXxBZbrPVR8arJAky0JGBmaNNQx5LmctAX+
hm7Nkix0urOAKuFcbHq7yX7FPvQXuw0p48F/5nuxdZOdo3ESzCTjUakjN9PPBuqMH4rw5ngA8RWD
cocIW0pdNuaeB4yc/9flxTxyG7qcozUhK4TfYX3rMfejqibBH1Aff4ZKgBnvkopqaImClThxJ7CL
eI+dKSCHnxwln44eSIZcGAE8+5yzIlM2Sbz7/wsZBKBFVrxlJRo/pMUCszaaio528wMPu4b1pE4v
Fjmoa1BDpj+FqT6Nc+hrRSshONRql9yiPCu0XXmqc+getXlsVs9jweM3bkKLmSWEJZXDD7BBnWyj
430RNDJdJbrwtegaJSUKT4kV1XLzRhQ+Aoymjj6CsG0GEnkpxCOgXFdLadoPXgpcMhTpNuKeT1lP
Cv5KTDym+W1R/vtRVf0RZ8fOSXJAh39exVcYN9ZqLNl4KsaXGVqzZqvFNQN5YeSfa+DomqFjlWDL
CgBBMlTOKYb7Q0ipq/OdYzs4d9u+9o+k3iruU3C80RYVqA5TvtSdz6vpbFXqC4KiYmLMHw2hC4aA
j/Mb/v3AmvboYYTEFQdVuRMv9ohiwMJ3HhmOLpsIYEZ6IXSpwHfHZs2tJLLmfmC4qjyjxfjSGyLs
dbxWZw6Nka33FLV2m58WUtqUPcC5EuMZXbiviBWhLqoUcK7dz9mRWE7tLfWx0s8R66+dMoOXhX+d
RpBohJU+DEEoKLwnxTl4cZuY+YctKN2z1E1G8BPRZZoYri2iMQalS7M85g10Jz+geLmosWV6ngSm
cguvOQkJEIE46/qXYY1qiK6DHq3yA5QqD6jCMUn88XiGQakX1U4w56oee4BnfBzUJhakNvm3A90L
2QryEhcVsDeakmn2PvtRgAMIzgtT6J5q3MRn6vSqLwlwz0DdqB2y8iGQ32lCqUStgf84/IQhtgsA
F7S/97Kz2qqiYl4+34OyrSlQC7Kti/POUu+ABR88E3CQnJe3uALwvztsxe/OXhiRDPPzNweSb+wf
5EDAScphuE2OIu38eHLVE+9Q1orllsNQJ9CkLRBfiTQvN/J2ccESUwKUWNa9kL6hKWstdaCoJszO
1ScDqNIerBCcwYOKxDi8HC8r6q1Oe/qm7QS5TU0W0nLa88h6Sn3pQAkSG86kAd8VldBXulZk+UVN
6qbyQrsM+e5tX6dR4elEdGvv5hVJMZFvfyuEmvLpSi34nLJvl4aaZgG+QtvmlL+ggVP8ta9RMtEH
fJRTVOGldH4AtuchInykzHd+JSeJ5OekRkb03A41S4CHbKIfbvjS8fFN7Zv+ClmESUoe8qlxWHCx
A9UH52tomiaEykiVNegKzKu3YoSySVwawbYNyMM6VDWvUt68rTsCRjOy6/a/DedkAR7vnfgNp7bW
xDo1j+K+P5hCl/Llk+gIFXZWx2E0WieZ5ycJV/WuvioyRzdbh1hb3ZMTgbgoxcMMOCwEvxvVorF8
HURbjE0P21apXVJhMukhjV/yuZdP9g96H+jwHWaFtTOn+v/4dsFrEVKbPmmE+WUKFaHGAk3uvI2n
A/rCsAvCx9kPzAz+Xtdu+LiJvZX480Xm/vO+7j6Hv6lZJ2ZVgn6cWCsGSXUXgD4x2IXGjp1mZarH
GLPc642o6Q39UMS3d793orc9vwhP+Wf5traefB3Uy45L11FM6pETn+2RtdGkGz9lztpFi91lHm69
yg15pOlx2v5RkgMCsdHZ6OVQqrW/M1Ha58y9AXX31lzW4AJeZvy/uqM/bI9ei0+mp7QjqqEKBRFW
JQC0SoH7m3A2lyLHdf8Zd8pPOtEhRXrEC0GhkubIS4Te7hB7Vxtk0CF1TNKBPHgYg8WPzQSRGeE7
pWaTmVmqGAlj3+MZGynhHJqREpSkBFIevFT3azOB5M5iHAM2kBaJM0HbeOMM6rYoFSXX/huKYXO3
0nbzC505fYY22oFlDxYVwtUlDSN+9GW/C6vYgo26Vd1ZIByOVqwC/Mld07BNkUPbgoCVTQu49VJH
7yVmoqX6es/wjvsSMAIHtb0acsKfhPNpMtLDFJ9avRAIW/gy851g+ilAB9hLf4cwsX0ZGWa+0qUD
9uR5KcZQZgBpm2SSfViqCtuEoNvy3wrq5FnflLxHq4dCcmc18HrbC+0BITk5voWxIY0r8NyVRfMD
2jGju8ROE2aCyyIa72kssYE5Zp7DKg/H78+5NZ725JgRF2r8K23rgwgkLE3MPMIYrijYOpvHGu8s
LMFhpwI2SkjISnIh/NevoxH8j3CCMvM+/ALkBwHeXb91II/3tq5YC9OUiY4kmZgB8aE0dbghsNKM
VAAojcymIkS+kg/S7CKrfF5Lv97bWaNxUprHOB7AnWVT2tf6jR27eMAJhfBmLOWE/f+OQ9KUawJ2
3yHhzyeV9uTP8sOiTK3QCMi01AKu4MGNEjij60i7Bt3gX9fXmoUvKUP8uXyG/xJ7dnkUvqTmLtj3
U6ElNiiLGwKGGxbJwBcNPl9qHOrDLdCN0r9gCjLcjPMc1DfgGNgAeG0aqDfZjejw+8PlNOq3Jb1e
GlBpYni5UFd4YNLe3R8rxW4E8gOYGhqmQ+d6JORRav14XCeBDyhxiqXVvKbR5ASSL4O+yxDW5y24
RL/fvrkRIQbSCNDwD9RzmfXdD4MBZnZsQA2IzsWmk088NKvUwTncCH5TXHanBUDv6Z3x2zUIte6T
WDDzJgA8vFwNf/nn78OqA7Uo/VJkHJZkFrbWS9q8FSaNxbeJPQ3dFlGRLtgN8qmmYHb2kvWM0+qf
azCc6R0T4ePFL37vU9//axiQqCzOWHWAMYaWmM3L4vGEOcg41BcxaLzkeZ/B0wqe/CEGCyuCAO6H
5ukI5HGv7vOHR+jm9mnnsk+rxKwZoMfLwH9uhONdzUG0pYsvtpj5o4XOHI4nxKvWIetjScof03Qu
/QVBuAGaw2nosoZoktWkLh0VcQApVzqvlCycIcHo6Trln1SIJY5SoAQVzv4VZLV9g95BDNDhu+zz
5Gp0qZpdtDFyZZ16hq5Ye59oSOBnvKlP3DaKH6ynl9qk78pwbBj2aAR/GNAAaFbqhFvpkoOUsAuR
rvFgMEwIClyttaRGOEe3MYmfOnRaX8PEKCdPUHUIKmQMbEcCu2sjDOR09ufJ0RrHuSCxJdUaKlTp
nrMFIon/bNmq/FRyXmarhHTCDrDtepLbPz67N3HITmkUt8g84ALLSGOwIN2lRKX+BPR31JH5L6w0
t42sXSkLkXfJ/wZ0mP3T+8He56CCnEVD7Jbhm5bo/GUDmulkLwYE6eM+PDFyrkcorpHwH0/VpwCF
pPjWUKy/kFLEjV9AAqutVRRG424ZsBLhvgT9GrqAmQGxijSbzFizVAlqQi7wjfA4SKIdBXChWic0
LqdtFVjrd2q5o43Ih+VrTKQl8IhvLgHI6Sa7fBGPrCsmgdSE2apNovktAzHvKOp9ssSy0mI88SyE
s+QOWU8O7GhlQOAVlojEMzLhpcGnbYlogIR0aG+QdEMAEzubyD+iWrG3VZCT3JhOjHhPr44ERszP
rMor44gKVypSJc2D13CGJatkSF+kue0uuqorhvqkMpTt432tXoaKCOnVIjfYSTaTGvebG5bo8SKg
vp4UUmTrI10xMTDyvyOfUMU9zeGf6LjqG5m1OYfEtfzH73II5d3eHFZf5dZA+PieD88atz0beWCm
d1VRJDKW2DCYMv1TrVQfMctTabgZQiHjsxZI7OXrnkYGt2SVimDCKx+j54nemR3zN5hOD3PZijdJ
d6K8+EpgKX7pPfXjV+VwEU/HquHjwzEwSysotwxnRIpWZL5Iw5s2JMOzhWsol+n82auPsrsRsQ8/
Ap2x4qSNXRXyKlNe4rybjweAz9xeJVSuR8OiEBZqP2e4nmrChgEr9d6AZFuEduLcb3iAVsj4ZQ1N
mzaTXxoLHxgBCbYJjHVHG4B59UtI5+6EkdyynGWR34UFhYZTa90oby8MALJZK3wmdrRpR87YPUDs
XN/SXyj4jNu8iWM+LHf1FXaabSj7U9DFzFsV8M7IVuRY7K/cP48sdxD2XOqzUQWo6nig4JNDDuYK
OK+d5waVUIkTyHAcx22U425NFgkJXg5TvrnUGzeHtw7ji/xKDGQ3z82S5A+E/y0NCVDK2YbgLj1D
uxRPKPSZ2A1ANUXaoHo+9c5si+jAti1RHMsFAdEix1d2oxLOM8RXco3l+CaWFT2vAInVAQTLo2z+
rebWmQtg9ns7gPdLvFoa03n4i8+G3f0PTw7+EbI6vKJffKLOO3oA7XPBv/y0V4CQ+MFtqpP5Ewy/
5/WXNHwphdI1iiEzL8HBG5HRPiZlFmgLfpSIZ8Y+1BOMwuSh95bvlKwhSZ8fpv1tVUFM7caQnZ5Z
hG8ps+LltNQjixuWokfb4bAGESU6/KEFerp1vyxAD4fQ8sT4h9ydDbKIfkZuxtalVM9pBxwck1Ga
5xuzXMcoPaFgDXNoq0a0qZN/R0K539D3pQASNETRLdT3VW7rmprmteGfmRT6syBXd+tNoNylRCLN
TfTtIAPIhj5SMSwuXmUtd/stTA81OAJSI+KTptwMI76Yv0jkcRMOWJPuJrpFnvwfKz6LCWKUnKvD
AWz4CSRv4FfubsRPHdSXDJFkQfHkiuQ7/Qs73odwYPJ19O31tO84OsY4+OOiRCvE4SFY04O54Dme
T4LRAxdoWmzy7pgK6jWDcQoG6zbNzBnbpd7MiEOMKfQ3stU7aVz5gXUb4Xr986/SUJ8bLwZHxo8i
9JivmB5gA+aHMhZPeEgrwY2OXuDbZYsNZUhPl/cKew1D0ldqgiDL/9y8Ova01yh+9S5orB/bsTt7
SFh00Hdqw5JD+1N2OgsvPgAy9BwXADJC4JMgHcKsBwu7wzwDMEDB/WIGp7JnoGdVba+9D5BZx+Hn
t/iFwyCgg9AZ7QBikRnXaB31zNAf6/fluS39oeqjDz49ZmgajDFdSMAIRBcrw6SIylfeWdUhlHeY
fGX9HZ0yYb/mMdnabsksn5xPSq1WBiKgWhagnBbmfv4XJFig4WrQ5KU43Lgs2+isy8wIwA72/j/3
uvms7d63MVa+JZ+ALuXjLrVNuBLKMdVDj9I9kP5YLVXNnEigq8ESgl7jPEq1wxPkY7uMLwLasz9e
b3/hL/tGp9YFvPEsePgGY58EelJqBivSNThQhBNr+ZnGXr4+C3b5dcBHW1HcYDGXEnuw0krTNHU+
zfUPf1EGEml8910/B616mBAvi4N2L4ZbOhNpSOA02s4qjfbu63SC+H45pKFma4qk4L4mCF3UEwPZ
O+tRFF8KwC6EpDAHTSv5SlvDdIJ4sIvqyLjX5HJakrcViYh9Y55/e4vpBo/EZ4qmw7tNZbz32/MH
6QTaquM1wfaH1lipjg4iik9HW+lOlFxkWpv2t2JKFLs1SyqZWRtn6iKzJn6OkEoHeaO6qODYtUot
M9iywZeVxWEMwjciBqXFnglq5RwjlU1uJFT1NurRVPEs4lj3Q8HkidwA9SS7qsF0XMYOiZE086XR
uMvhNqIFNHVu16CkzYSakdFg37bTq+J/dfJlEoniRi1orgYRdB6zyG/rZfWIXCQenrP4aIgMlMYz
SWlIAicW9rmVh5PFkAeZO5z4BKXvgninTY1sl/w0WR8s8YO+vZEq3CL68Re1/zX1KAXyfxrNgN/1
uMd8m1B4namDIFxibkv6GOq7ClY86I5p61HlpaMrJsbcby6gYH7oDkswxuDekjpeiuDrGoSsvBLO
hfGuirm425Kn3/dkYP8dsZTgQLbEAUvEN6zTTj2L8POVcnW7I9ZX8QOB5zGJvU5lhmd0H3vSezqd
XV+Qrg5E+/BjZ+TyRUhvbBCuCUBTFIEh+i5jB7eZpzQ3L3q/tLL1ZUfKz97xVNtfTfFnw+u9BS8S
NhEIVdawd5Zw7PssPak0xtIrWe8RDrmgQ9WxLmdFFIzNX1LiGYwXbs8Njq9jhnJO+esD24bIUNfU
ZOQ1p9SdQpmB+YCXsHfgox+E4sXq3urkbAwoOyaZoFOn24E+ngU/7jCxSCIoEHINqXw7za245toE
PUhY9sgT5gdxFyokVXRinVsMwXTi7nTR3fQiUcRWiTLhcxRp8Kgj7JSQf3w6DmT6ZZwEZiip+l//
9NtKkMOKIii088AwJTc78Gx5eqZz2W/PyxEQZiSCkp+85N0CWy1UZoRoWKOrcIscIrGcFofT7Nf9
wXPEvLBMGzxG+c/G1UqE5hCFS6QbXIPf3fhCQbDGzufFJRKw60Z0aiYJzVwoLmB5zksWHoQVpO6U
Dv14o+yrdNVWZFfZJtsFL/C6D4MPEg4LSQIa8hJwMxCerx8AK+c3BO+oZHTZJIFwpHaUTiTYRRO2
kzwkSWInGRAaf/kW3HrDBifttuIWMW5gpr9kS/rjfBIIgdbd5UQq4FMMuCS0ZFOJkbLv7mwSA9Q8
v8Dr0PjI1FvovKB5q864D88/W1k5fQmD2RglMAwlcHSmfWdbj8n2PC59lbFomv/WaPm94MQ0FXM3
IP+tybvMx++yn6mDtK/Q0xzX6MW7Dn/PqWmXRi/kdBW3gE8VlJKWJX1EwYAPWZv01XxnCMtFGEtI
+NuCGTJM3uYMg1A0SQmUWKiD3PJTOqvp4wtG4T3LXZr74chVcQuSzxe2b/ZrE5GC7Ik7sTsEOVPd
g6UGID6pvwlvLZ85181kvM0UjbqCs/CPguRkasfFQ1vTuB8HRpQVA8W2eoJ/ia122VDd9rI22yKg
Qv9xW0IObAMe4v7/mMX5NhBmTyMpe9MD6De+sM5HlX0Ft226yew2QLRkB9jAR8bQBeIZ16oVmv1F
aewl6xeh/LHKTkCMB0p+CuhtSXhl1Si0ax3qrjEpCeKjfLDV58WMI22ymgpcMrSbn6rFTwvFkY9h
9h0VKPEwtsRbrRHAX4YSM1NlKd2/sNc9xBjhpr0WlPMJnRv80WL6ofuFw3PIbRd6GZLybhxYARZw
5lSVltclkxaIDeE/hZLS6HQWhvMH3FYAVOFdQacYYf0O7ZcYHG75HPjgwvG0rN+zk/ExtEmoWFsW
04Z3nBZ+rkzGjXBmtqgW164A6dFM/oGd8k0YoyftoMxVzRneLEoycpjAbimixdBY9IiB00izRzs1
wrE0RcW/JE1qRmaQ9dKP2hhnFxQjdGaI0Un+kc8lcLzn8Rhk+zuUp8mS9LZ/SfSFF6V33wc++Pv3
v9aZ0Gt3pkhLYmlEVj1tr+8WQMDMxkrKF3JkJqtesYjvBleH49HegzNoRLL8fDGukaOQmUwbFlZ9
h1mRrBytCDNhq6oYypYnYoDnttlMRpGZQak99yQqfJ12ktccLsTbtTTUscu2tiqrVNuKydjcOp5R
yf0fkwfm56Y+nQZKtMEhaQaDZa83ylnp8Wo0E8H9+mxQhiH+17vNUQF9y9TsGuE6URYhy/fr5wiE
H7vf7YP8NjDUKbhspHu3zSPXsk5BFE62hOrwSZF7zsTDqcQ7FJRgHGlo1k0Wxky0sNTz/aVsovPN
l9c8pTawHVH5qxMzw9+ZMH6t4Fe9dBQmqADwW5DHm7FBLKC92ZKi9Nk2ZeyTdcDGDMcC7wTGF/fq
fD4XZVXuauIXddGsUeHA8XGiVLfOyOElpyIodzNFiLaN+skfy4ojFk2LEqLnMXQhWmO4VvkMPAjF
HXYb3ipS97/D5yvyN9EQRpqRwJSRtF6CzOd6aZop21jQjp8jD/m/IkQI6w7TeOm6H61Df6AvH2Du
4y+vXMaRKwkgewz7FQrcotRIACvFbq2NqDWccuflAcguAUTaAoAdepkroYNQRQZ7NNpkSDEQOPSX
YoBNdoR+ki8KZkMouOHki6YnqERbaghOpsnMA+hi+eGDBoSA0x0VeeE9ua4nu41OSPsNtwWxdohw
NMAw0sANALdPKtrix5Fz0KNyHfXyHSc7Z/q2trrHzDCTBrfADrCO5NUr1XDR9OI3PDLdoJPOPoth
14zN/q+tFF0J1H3amRMS6Asv/cXYsRjuhlA1tmnCeosn4wzN0dH4ZBsDhqweq2DOFPv17pgj7Wn2
CZ8GKXyaQ5utobN+VHBsZbQqEGdaq79V4MpTfAp77cVQNZf76lFVtik5IrNgs0s+lzrutZqTMgZh
K6/UX32cesjDRs0kRuxBWmd1wPMy1BI1GmohUm7lpYxcOMUfdj8ZzteuP3XeVOLs0fkBWXqjOAd8
BImgxeOOBWUt6tnli9RF1A9Qua64sVZd+MAIHNcNPHrQ7Bzhr3gEZAQHjPua6OoltbiAv9GuTZNz
vvgoXahyfIoOGK4hcOlTEfKIAxnqXc1yx+nbkilGCBHmrQ9+7aV+uiXDqDpFLR2YeLU8Yo4sJvzk
3SD7Op+JWkYUXliejBzLvJBUGfmd/eOxkRqDPA0TKv1erI2N/gSIVrsHBSLWH+KI3NQT36WXqAkE
eO6Gdg5CEtlI96aAzZJ5VAZ/HEEGZ0oRQMfGrf9PKI1UV7JSpYSxX3LncbeqE0OyMMJi0R0aD92y
6UIQ59CYJZhUkiViVLesKUM8KnYgwoZp1Fw7VilNUD0nwaRQ9BOAelhXWDNYDdz3PMyJRSt4xD09
pBRwTK439LrhrOW/5UtNluxkepThMn3IePOpj6D4Qmhn1q/iHq3VVfVXySAcBLTn/N+2oYDnQkSp
bFZGfiPxXAFv6pubrfuN+gTnuB/+DpEi4ir81Idl4084hqHLc+Qdl2wJmy09HHyzkErEYKbrzNTu
fnbj/bCoIbPFqoubYnDvkFs8vkA8fvhcEbJmVkznGGyBlDQVAXKLBqsMDOcGo3QtKkO8sjPbr08a
3D5WyVeSdvEBHOeecBmB59yvSGnfZbVkrt8IKz9x9ZmEiuUfq7gPdDAJvmmh2/UUH4zRSOhI3MB7
cmNqE8KVwfIQvUGjSbdLPJDqxV/L+VWnyN3ApKWRplpZGto56LrddjoptPTholwUbcur1lKwTnf7
q3qFiuX1XhM+fa8eag9V5TTH0Gd2j7SZycfOSzzzGD9PAzdnm5Edi0FXJJrtRLZmro8rxienfhtR
vYqYae3JTreDEHxRopCOOCOeUPxEo+3QQZyooQKl25rtmFDWAmGj7yHCAolj+681jucwkWDKkE5F
bqFdDhAVIchfms3L95bvT2PpFYc9X+rAQ32fJs1pghPK7+xKn+zAHV+hAEjhP/4Q6wNiKIBgOJ/D
LidoZtozRqwfyBv34z4bKJSFoYJ9Fkvu3+1Zhc9fV43tA3Jegz3oEO0/XLRga/+F5WW4fAYkjNa2
5euPaGWKiJPTX65VytbYyS6b2Yd3Wkmlco2Rp8l+NjIX28Z++KFi2Yml3TPhYTGwrUEQlteiPj4f
uhvSrMCUGwaSmgRZjEEoRLiQUO1WqlTx+Mtf+L8A0hwxxc9PzD38ekRQvNSKjzIjQOkYamo0+xKY
owgmFt9VimlW/M7oB2yQa9uGkY2xCuE3wO3OLAB8JZCyVFrthBvJ2lxbanRtXSmoAkat/VTYojeT
fusffJU/NsML3YBPUokIf7OpnmxyWHlXrWXmZQsN9eZRg/DXaMdU4FJZMabx+Xr/m53aV9jjd3J0
j7j+wFUjx2lTA7zfT8TQIaZkDRH64oeMSvL7oP+lBY9eE3bcgs9QDOP0MxP+PDtFHXRsiXEpt3+M
kHPUNm3thpB/hztxqx/7We7hFi/pO4gP7RV43dNxuCiQSBqgxj4j7SWFhSCjx0nUUUZuS9SYeWgX
KI3o65tkx7kB16rYJBvlfqesXr4cQDqOgL12ddE7WlDRIwhl1XwCW11IeLMA1frM2g+xEsaCdNTZ
BxZMro03EOqgjPj9oHR8vTrr4U+EbTfV6EXWdO+NdMVWa5ibajV7JEPSvBzG++eGMIFHOzvUzOqs
7BGBiswEMz2jL9N8VgHQoVsSI7xrUZ/SedfMhNvTGyzDcjJ+kLWbZgmE+TAWB4qL+bbeoQRkHJTu
qTGI0cbY5U4XsKMFjfDG3q9YgteyAKv9d6G/Tvqpfd4afc0zbI3Bceidayb7yAEP3bvF2jeD8q1r
TRvwfU4QRlN+i7QldKwcNgLSaY43X0fkv6JD35oAy8eF+qBI81kiagwVF+ImO4lOOfpxRQBGHKk5
5NJf8iXQP4+4Zsz3P+EzDjft6OByKEjOACnrlJ/jhBfev9Nz2Y1OM6w4m8sY1so8+/f3OAHPmYmk
m23q4tUr4/1XRuH1CW/oZnDc/d7Vvv1HPT54H/qBZHjb97Nzd4jDej41a5H7crRulWrnoDalwGKG
380MIK5DvsvVfgMKku+o5/WZ5/w6IWmnyd+GeCstyse3stcf/sfVpNZVIwwLrlRWn8Xmw1QPxMLF
N9bpmBvK3dMJKIt54z2NObCoLIZE+suDdOp+sMfhTMuAyZkPTfurNy2S9vZv+RztzS21tmq/BxBQ
gEO4qwMbNCFixxV5YzfgqQRvqPS6ePdb8+lLAVIiS5VHkOYkRbB1U3dbGn8WrrCakDvPjVTA5smg
lSGieD2W3cOjC+77Kkik4Phzs44LqPwUq9+RLiS4NMsAAvl+SdS6D5IHxDujQe21mOB21CZqxyiA
o/hA/Q6LwzhgCzAMrViGrhCri+75XX4N4Kcym7KjygRk+AZ8kJ3xUHk4gMG4y8fvCbSHcgt3NcZF
TuFh0H0fLfrky+A9zSffDdR+wnek8ZkovR3sMMTPkMMtuQ+JDOQGvOCq4v5vUMrF2Kwc0eV9c+td
Fhip7Y1vHaEEyTRHIYBunYfeWB4Fn8ZuLgWuSJ5cIqJ6mFAIghXhDUloLlm3hD2BzGMq/wKJpJvA
cC1GsbPc2OJYIrk/wqdhvA8iNyR0eUTBYeVl3pXCVmOBUbzPxllgMGyvGwW6Yky8oNcw/zOEsKuu
CXGjoCXHhtVUuCBAebj3ytiQeC5ADNmPMLLonW4n1xhQe9zbbnZtVwBJYQxMzAkciaD4NcUX4l0t
5PK8AXQ64OSUT1nXo5J0dqCjGsvZiewJtXyHXNhXmLgI8mbeg7ceZwV83/C+3NEPLdTFk5AmpMo6
wiEcyFp6znlNayeL8+zZPJhtvOzeogIyVo6+se4hLQTsW59QRpDT7ZCLCj7FcWPy/QYpG4AatQsl
UcoG4Ubtadmw6PXNvYq3/TlQLh5Mef0V3a/2LYAjnSdEgFMhZXjjJpy+RAWhsWJ8M55wV9wUg1eQ
fMVGulzZ9INZIdsTpaU5lDHj9m6U14++jDVX/u7xv3bYOttUMLVrHWCVF9kOfOFLUgSnEiulxY2T
hZJCp7Us1TQvYyAoCc5oyhoOSPEqukIXSNSsV0x3WXc3a00NKIA8Ehc6iUHog2IdMZ8aD/FMqkNw
fCa0+p+BrXTyhu3GrQbYro+f7F4aXiGYB5sAPVz+CB724CuRTfF/ZBRL2idN2DD9NKfCoaaUNFet
R4/4zK3PUjiYOPrTRJP1jGwRg+LdTJmSWFQCSJX95oj0G4wL4d7mA3sK1RYUSnXIJiYPgh3tohAO
XKc6xdgnzOH4jZ//2mKcJmfR5st9h3sla9UMsioE5RtdMnqXfqDP2cAG31D8+GZRt/i39JZtVDZq
fPSR6eMtnYse1HyujdYVwc0mWaRj322szRFORGywXbjWGGjLJUFTetq1rqflUxcDjbi6eXnpqfFG
f8lo1rPVUQ0vrT+dNk/H6vin/QBa1LTVpVZ9Td57hrGeatStVMGop6h/25GO5IDEMAAycdradvbD
BiYSqMXGtKWXzPjMLXW/pNCFVbutJDsqij3eCMeFweVmNd/iFFvE05Vd2wswfnLpNDfwx83vcqeT
0D72gXzJEuXy++WiTVz6wSxaf9xeAQnZE+k6ey+wrIW779nLtKBGj9weQQUQ74Nr34NiAnFgFzOb
srZDAu+yusHpJhVa3277jUdSiOGQIYAyBJMvpUbsv0iefYSY8vqOkMMEk/UKl5FYD0Al4EUzdXuC
fQ0mIdp5HDgSpf86XskRdYJ6QU0OdSHfiquzVUamVcc1BrvBNtLwOQiX+gOuXRGwfFblW1TUZNt0
8MG+geG9sQs9kB1uQWM27kg5zutIRkEpZMzVtdAjl2vTRfD9qs9Wl9yVKXJXDH6n3UWsS9SfJ2Li
RLTDaNlqVYUA5+Ob35YmbCcAsxxAxMvyF2TzlkEw2QL1wU80L0da8DfhmnvBAiyBm4dgr1V8a4aJ
WdyMzArZ+evOlvM+AuKvRtbZph1Sx00Of4CgGTLUdnsVVLHi0qD2yDJAGIq95aEZM8dGhnJotToQ
oksjKJT+HKUCjOXpX4KMBhzVvDLrdMgc/nsRPXzA7zHjnH7P8vievhFpsDbUv9s8U8/GEMbtGj/n
H6EPJsJvi4CxpE8z7Fyiv58cD1hthOpVxdfyMUFK2XMUzS3Tl1E9Ae5WzzyAAnCVKFCFZzoV7mdU
kVrv0tfP7zt1o83DmcUtlbszc6TXtJtFbOekezPvS5Yt1PmsHZvllzMyWGz7IWh7QNUNARdPOSiU
2Nh5DcLWUVuEb+eEvYGkka1UhgYvsQJh/86kRSTEOQGb60cRCijMJV8zK5tS7cJFpnw+KrLSOd7L
sjTC2QMLYlrle4NWffctc0vIl/sFDY0fFPyr8vJPANcycL0AaMJAB3Kdl7br6KjtDXUPlPdrk0Y0
YxNqXXsIHlJKgPgXwpXVLAcRzqJ+TOuplZQ8nNJu+h8cndMt7Lpi1T2cL5YL0OgMiG6WaaoO59kK
JinOM95vOWLnHXmw6aGJj5dv8g1n/e/9k7M5X4owqPdubbPe/EdgRQMGd07T0LsihXcUXJaAoDy/
lS5JUbRrdaNI9yQgltQZWFiOuXCEJkyNjY40ohRM96I1kicz98rGUptA2yztx8pynJGLgDTT3f+o
beizZEfnkhYZGL+wsFK7q3nVwiuHf+CvWs53HRFz1UGteHdpPs6h62xkdamVmAb304dwv/aULyNZ
srgoZFf2nS3Qt/insfm4PRFkmeQxLnKCK1c9MQmOheODe9UdnsZ/ogI69AerQpA7c7ItpbA0ugo8
a/IO/FOX4l/PNYlSllhhrR1kh6Ue90e7abVivgGvybBJOoiz84NDzZJ/+CQY3T5o9eh0HAePAT6m
79vzj8+inIBJNt1PeK/69Zl+VF6rfZDdwYcrEYR8T/SvOLC7nCtE4yKFQ2G/tlmyP3LEFrTfGcqv
CvyjzuOsnhfsXVCKlr2c7NAtO7nbc0oG5Jz5kYzilQrUMXZNxnotL9faoMD7a0J7rRtjDB9/WSKq
zNWAwKJtT0wE0yGOZsRs7ZJIMUHGKeoLTT8vgwA4y8e43k6Ckn40U0bjBXE5p5aFCceEq8bp1a0U
YmPl2wy21sIWm925r0UTbJOgRSmKY+16bOZQXbc5ZLDj4CqH46d7YAeDZvnCF7CDHrcl/kL7vq0Z
aT36T0m0Gckm8fOwhVDYeNt1ekGWbj2andXyGkAu/XMbrwdKFCU0m0LKyMwtevaJlrTCCxxYc4Cv
+/1NMoyQkFQg0UZSsLCYD3e18OQR5AT8AQsGoQ0uW+kQDxJ++QEhOmA14IXZTDXNdZbemZNmvweN
CHKC3v/XYfwYx6TeUcAV72khk6azJTQnOLIYfnAdYIDPT2RkNNccQuhr+XlKpyiBSGtzsb58LIIw
SJwVgPu9L1JFoOop9IVXyApFglN73/eIObmQ4vU3x9yuKdJnx9eK09QgMiuYprPb+s+7T6X8dORp
yV8It0PKYYjt/YTLhdzG5SgEXjgskReoIuN+zeUVqh5jykNKKi9fbde5tMx1qHYPz2yj1JyHF0zS
BhD9mTV8Xqz9EkWKxzKPoESk+VAftzLxub6peUhMBS4EOsvFko0a2j5fBM5sv4CpoJreM5ASxnsf
U5pmKIwFni2mvSl4y9Ry2/Xt2MQyjhYf2H9EHxRUeL2mvkElOGbNfnzuovwM1r0HLWYBowyZWfPC
67jUVXqMnKtp87zfpJ28+aXMqzpZpBhh8zJWtabf0zKL2WQnNbsskeIOlL3UPRsc324mmAKx424a
iq6D4O0RGLOlIhYAbGVRhx0Si2bqyXtBToP3V1tWPTw9UqwLgkqGWetwZnolmHeIDsiLTyxtbGjS
Dn1gKer47SxTbxeH5jcY/PDqbBvheiDcpBSm8zydCfMi2nA6bQBM7OacNyhlg2xxIw+GXGueUY4N
WxyGa8t2QZXT4KMNuNxN4fYwDjiUCfJwFPeTz3CfXvmWXmxKaqkWZPIqSd7pNKfMNEYPkN/U8ltO
5LGKi2l2evwey4zrPLfYEMtQp9yx25crBoiswKDe8re5ov8T5uWXwFLr4XNfIyCTStAXoj9qMrpW
E8YEfukxNpSkBFs3v6Lz59z2PBJ8mwHOLEWMizCfaOJJo5wAkoyYAXqH6vm4vJcfoKhl5RsD/u7B
VMvX71XTHW3Xb0ZicVIY4eWyhE2zUCXGhSWy2JJAF8wMIcg154/2m4QWVF0z8AaqlMhLJ12P94Kz
60ok3TGDsQNnHVzA37p15sed0SvIyR1ma9KZBm3rSiPvxjv4SQhB3IvgIwk72Y655NeeDTGI+I1s
60/zQfsa0dBqTCuZnfZMnZS5QQ+QIQyqUeawo9wLl6Bfx6uOFNbk8R+YMoT7nTcqj8zb7Dxj+J0Y
FM8pGBoA7c9Xaf7NSN2LjpX0lMEyIy9dzayvvCa+RE8sFl1o2b4bqaLfQqB7ysPf6jhX0hgTWOmJ
fzgAkBXq9ROuwiwaHP2r3SPemvq4qDXPYihXisVyfT4Ul5O8pWxEc5tEQUbM91Pc/4GfvAhhRkhG
LbHDfxfEFKhMukKYsXELcxilM5BKN1LK9pySv4wn2yIqoQnXjJh8gfqnygdFwW8IM+b5E7KYGzHN
ILBrgvCbllg09XZvof6rIkkB1usuFz92IQN6BSCYsVVSJ5VpVunMQlcVPn82MkXs5QPB4DNuox1Q
Q1hrMyiRoGl3XngmZFx7beZziuIi55tGiMNw0hluu88tzIcNFBADl+rB2DUnjbLLsswjljwx2emg
5ht2RARzxs/WfsIhuaM9vHDZZEzmiU+v+6sgi70X8BhTkqFbughMleU33w56LTM3vkI+ljqvxDVk
eJydOovpuipzVuG7vkwKzZ3Dy+btN2u76E6Md96h89TOH6txpWZIG7puaG5F//IXrCP9Hkz1kPDt
ADtLobdJnYuryoHmTJrzJbGCa9sFHnAkgtgPev0d8DG2ncccXAJ1bZVgg1/w/qKrJ0PHnYqdViOo
QdXl+MuI79Cm2iqNG1dEZLanMyBEv5PeLSQ29zZRXwqGakr2Pf1+SY5knVWB1VpPNkk07DjJDjjQ
VnhBNUMsZKMB0k9eILdwGfMZWNJMZ9zwYBRPT5fSf+KQTDUkH0vEdihOQQizz/UCDW73ipkK4DHF
LSKeFS9rIt3B9LibCCdFIcygc7Z9A4gsLtIMcLqfzEoWcwwwGNN3KdzQf5iz+EStvuOxozBXb02u
/8FwX5shcDEU+tOkrZ9WuJDRRtG5rDii1XqYVyCsmTu4K9NDCrpKetWOCBohCpKOK7l/aKP4YDcd
HpveqfdS5zlM1Vjv01g/zfzNZtyI6ut7C84SpxB1GjfXuXbUggvABlTvA4yg0l2GD+htPARX+R6B
4nFhXw7ZOI/HKyUMQggf0cKCh9G9kAr7vECI3is85Zo3J7eMEQgkZEpVUSoVwQaWOsolgYxS/hK7
IQ7ZH5QUIpkqBbXX7TsejqkaOzcRr9ILvfXzHoxyQ/1FHHhHC0NxYi98+m1O3AuqNM6cXw4ZpDsd
yMMptiK++4nE69pWjn0OTnQg1r+E+C2AvvLkvSh82ZrIn/fz8h6hzg+P6zYl3FvTjnk8W8tpRCC3
nvH1Y/nWjMGttYNr1ixLzoHEHo+tjBU9s4z2wJ8uxaB53Cp8Qaagc8BQMNkC+NeIOVoQHLjp18Du
hedgZa+jlon27x4BrwNOWa8opEnGuei9am+Itad0ZCwFdc9RCbLp5fo72Td0jRzbXxIDRyj8gtMh
YpQvHT2tBkW+CpRASgKTczosdKj0AhgP5e8HIUCUwLZkvPRbo4oq+dcaf8vbpCfsuWLG9wFAfAQ7
x1VwCn9mlk9KiRLPVlmuHf73rmjFAYfmU1hakHvmRzT7FT/Us5jillf/w47BRyNBhxtiSsScvCvs
torKSnPQheOTAjzo1NcLzDEqY8LHJuGjTHB4xIqrYu++N8GXuk3uHfuUHJyTNLsJrlNFlcr9DmI1
4/bQXQ+VDmHTg3HaYmhzYBDBEucv0qcP74H1yzeQG7XRhP8R5L09/fBzJGQoh73WH4FQvn5fW2ih
U2vWbB4mxKcNtNJDJmEn0KM0z+P9zbOYIqeawgTzcqVHNeQjSfpQ9eqUuhLgFDfkxYToU5nL1t6J
4VI98nckc3SbzLVtqCH0HXmWPFjmQBDU+pjIClWU2Gn7dgI7aO02Ohfg6SY7/Ty0Rg08CjgK6dlt
T4yFQGSg35oNGmH/Kx5O0xZzV4NXgUZObxqO+oVJ8mn7LdXaO3QsMKEj8jryfUj4aOPhvBpHFct3
B9Eh2rMVwT4y0CHDHn8zYDA2ObnCHG2+ajpSqiyVdNdXvP2pDq/Yf2UwCoQQEIYYwrpcpcQ6a8vG
6qgSDMepZtkNwC4NdTE/agEXJCuY0cuKhpVAWJ3bktx6roq96sBSdTONxv43us6A4JRtCnlYUtLE
N3LHrvWRqEqf0zyp25N8WJ56wdlGfEAI6b53us1yBCNR7jL1BYF0CXYYBfTxPEaRM0jvuxL/hAC+
j400XmZHLLX0LsIJDoJ9sMG0sO1idM04oEdR7mkl5lrUj1Rgd4fNhr6qAOwhhv+LG0SI2goC9C+j
3bl4jjnm4YB7TFbOu3s7wydiVsXZFMRqslCUWE9BT1WdxnBsniCJwVxsb3T6gyjwbGGJ/UL/hhLw
qhe8REPyAbzTTwluQST/NgMAAX1lHKAIZizy7RSJ2nRO4OKozzh4d54XepCmydaYfpWdXhkU7rMe
c8KyIU04qDE3frWz2woVlhT8u4NgneuhcTgTWjboEoxVs0PlWe0M8Wk2NGrhCW/TM6f/sZyJZoer
DXkN8gZ+TC+ZusK99zsXoU73fthWx+wf5lQC3L8JrrbDbQIDsOG61Z2wizdHpytrhGEO9AyZ35/D
bB14uHLO8ewduGGbf1wzLE1ZnJZec9Ele5jmDFez0Kc+AG2dw21M7zht+J+3W5LLJBpyw/A4K8+s
d+DFJ8g+JyDs7VISG5eA9qEbUdlNodvJfBoIox7+b9hDzbvYpZG+TiwbArCrvNCYdNRl1L5s8zqk
nnaK5IPfUimv1UhLOvE1Z8VKrtoZ0YVxOcyhrM2WRs+KOYncrivXQvT9uxzZ0zK2nHwpk8Ed9WTs
qAlp3iQX0DM1xadDuj6r7pVgpyKT+TjhtTFGatkxzJS8Ru0HfbUDP8mEOEGdenuqFIZHoG0ohn24
1WyzFcne11ec1dWcbpZQNqRySevhn4SoBiojLl09X6rA4KuezrFi6akBxAf9j3UFDTAbDkwDiVuc
JtK9lp9oZrxvy0iOEFmL8UNwjfJkl5z+RtoaSiEW7E0xsWvNNXyFRf7PWvvYZcGRemvQWHwfA5oN
B07HllTSnRB0py5/F7c/gydg2BFUAEPou4Qr259C/duKu7I2L5Nkbvd0Rm+pUOP2p2cYTQoxSMis
LBb3jqmkUa5fs3hjWyS+mXZmHNkE2CHt1yeSWwUWPD1XwAMJw8x4LHazUw92Xh9/GqoURO74zwAO
aUZF5f59hEQvCRkOfdufqatUlDHMEWHg1KZCVRwMBieO5Tf7S1UWzeKktTUHjdJfdJhtRMsKfaxA
WkC+3M3vDHICpML+WULV48Ut9/lqtxM+NfXvA1KnaKQTr422kzu9t5/kxXqL/KTImJD5qa30cwWy
JdyWb1VIMB56wsFjEgxWqeIIstc0mJvz7VIm08yhSSkwNL1NcAqR/9F2iXbs5r3Em4vrlZ0jky9K
J7SlHHfyEOaB7parKlj6sTRVz2oeKvrkWoyApVIcKXU6HtwFI089K8DsH7wdp6ay7WfVcAw3qhzx
yN6PvNkN6ldVFvVFSd6SqA6EUUdvfvw+u5Em8tIgVGgyDE2mIWIZufqHEj23OjP7EzSA8vc4Fe40
6lIheLFC4W3LTgY45WfJ10HWYRoKjF6SBQaxhaGHK+d1kXNRYxMsBZ7FNHLOr1u4XpZ0Y9IoeW06
R62Vx/dC7/7zymy8OND458z1gn0HZcTl4atpSjYBfg4he0PeAXLGhFnfzWsrw9zQNidQ4xYRlud8
PmenVd62YyXzz8scWRcE1/VqAVTokkuy2szOOTR2LyFd6fhLAwCQOV6AOaLA0Ux+O2cUf4ShkeV2
pDjv5aN0CHYbBMCbxRX7yFIhV9JzG1vAdnYvpzHdgaRazBpjeSgg3kJS8j5ox/fMY2Lampm1Sm1y
8yuB/SjxV0vspiXS/8ksSpH9+yVZVenN0KvedLg1d6GmYSbe949LjPue6F4aBVoi8WP8MJXenyH9
+1w+NmXgeflJYQQV7N/MeT2rgwViwdUE8lTJtD/ztXz8RLC9IorZhazW0cKkV0XKfrQdqcKMPTrf
X9N3eWG6uy1OvDjJgi96AmJjXm62GMxAlSpe0Ek1PXTYj3t6hqYlyeTCZR9QCMbcN3DSucIC6G2D
ckUZLAe7zxb9zjz2Wca16Hf9JgeW0xK8LTuhIWiPLn9wrXrO8JMhtpbEDKOiYbQwbvOQ90HqY8xn
9AfJZsS5d6o+zMeX5ql3awA3aE2wylAX2t39jC0KxlSYdQeMyDjDGnFbE8KawolX1jb631EBLrh4
6ZUlz+TspBXmfMhnwnCFJE4UQQt26mZYAqQqA5/BgfhO/lkKIhSlmYw9asuoGNXQKTasGEEb2JHM
izd9n+CDMij49Ble7BICkcnuFG9yfwj8XeIIx96b3XISsBsOd/rb3x7SGRywgJixKD+umy5oxEpF
TwvnCD8t/QsojKd2OL/UnmvLo2vbKOH6BjwDKT5AoWvFm/rNd6rTaRInDvicCYYStV99qb6gtIlE
m5IsywTa3n5otb0nSE7AyZUY19XoNQHF+a6yzp73sx+/tbW0mAo7BLXrAc+aEYE6ruTx1Gn4pKhZ
DKUk7NLzoNCrBTJYTAsmnhN4bKg5NOf9puESWhiQg+RnGKxbTK9wLXeDTo9eOE9UKRr6rwrOdT3P
nYHgsoxFK4pXpeSrIRNSpF3w5ktcoYx6+RSkFKQXlgNTXBnsZkkropTvRQQVQl4K7UypQP1w6vDf
f6d4JDRvQ8ZNPNbwvAy1/Mdg/AGXundomdNkwt5nPSStsmBpHjxCYzizLTHC1mPEIw/2mxsd9TZl
qn3d91SK8ZpWmR8gqqO7yXB8t8XgtFy92K+FXIK89PFmLO8ou3AD2dUnPHad9CXwGIkJpWcIU+FW
t7VM4XMVdcuTr0tDYujm2ltdkvS1G0izubXsxD2+j7Zp7RjN67BULJg1oHfMiyC2GHbceLTRRWU8
jM28S9rD0PX3iMqrwzuZ8OBXeCEMth54AexTj1FtX4apX8wPniKLcjSV5y12M4s08sOUsNTT2+k5
IMdrfGl6iLhwSIfvML6+rg96e5rJ0DIWWYBQg9A/inG5fFVemZbelhlwVuaeJKqUURpZ11iWtvNo
58TfIFRR8peuQshrjSkkx6kTZZ0Ox+sjSXq1UqVocgWiEABKLQ1Mk7d0aam8lNx4zjm6Vo6lW8oB
T6Gu0JGW1O6Yc6efthSt18SCqiYxTvJXxrfyqI12LcjoA4uhQyPvwG8KcprXV/scJQkxwT1tECLD
8ZEHBERxnwF5VtXEuSKDVOzn/JfEOLGaw1xFDIz1JPM6pT/HNtMyBx5+jG61RojCfPxMTQLogwH+
DwQN2s3Cikcb5gmRQnWE99257NReQEP4CU7aLe50ZEUwTsDGb4H9q7i/iz5vYLyfR/LgB1Cwhvkx
yXM24ZbsjcSyLX602X5K6D7cmIr/i0zOI5SVBaE+0mmz69hSsUL00ZZniAA/ILL/IvYNp4iRFQWQ
7qphGTq4c7wx/P+y/nAOa7KYdHLyP44PWaFiLMRAN6N/SFXy51VEFk3RwDKeImcj9gNCFOTsgO03
hdk0uJ3lYDx2Ffl5dHrchGtoRgm8ni4fTvqkNJwZGhkVZLJpzG1XwKNULKMXpa+orvj4eK2hUakM
mf6wkhiWKddTokWbYBK9dPZi83ruOYPjmNgxUMZMIuFlTmfkXI38PeK4K7s2vp5mlZBpsIaAjwNr
BUkMgPMzQU6KAHi95Bwwo2ajeNzyVr26r/ruySrIHRSDMVqW+wWk5Bk6HoRFzXcf5WIl6WI2tCV2
9MCR+keeNXCzjCeP8215YdKcW+NihzStJ1Otf8hzx3sqG2bHkHt8sqEfw5L76irAMR+GS2tWVZlL
/y4xBQaPQ3JzFsF8QwcC8RkqlBjmE7L5he3aIsE68g6spEdlL0M+gTmJvRlBUb0hbdYXEJL9/80p
CFKl9T1wf51rNY15HabQAAfkX0rjnc9TxDM+LVELFjlUicWkN8KV/6aQozVgW+7pnlR23Ilcwa9V
aKec3SsLsDQgkH5X63qcAw8pFEMdIeXYKOowvZfn559gkuX8hhcwX1tO9d/GP/2rGNI4a7Y1em7X
Xi2vJ6ivo5E7kagqEJ0zGOFTdEhaQf11e/VUfdnzn9f7hD+dJMW5Ib+90DkOwX1RtLqCl0ZOdFtN
Xoj2J8xl2i5Zox+cER1VzEsB8DFRi0y9/6AjZPG1mKLiD+KzsQXjsl1IbCl2Vccnp9J+gPJHNcNz
1QvxDvzNHThvTwRyDpjc8WDQvaTkhW7jBeIKOUcXOdU6jewo/Sj8BD/K40wAvrHJp7WYVxapP9nx
QV5BKg5VAhT3Y8WrUwSPJ5cmHv5xGKps3haWo8ibdH37oWkuzscaYDnzLPo7q5IhINFWvDeLFQHF
4VJ3/664mpnmlvcXnBH/1PBHB4Zr+xSdo+ZEAlVp4mPvDRG5MYynizpgbBK5pw5dwaMlvEWKeYmP
Zdro3JyP9PqJInEH4q6LSkAlpP/olaUy44P608oRPaASI1lMGPIHwVNkv1gKcjyxzsu1IcLy16Q9
9GVL4mTEmNRbMK28t2da4/tCrvE7ujQh3X0jV2Tyx32c0IwQkq9w+Ra3stBqZBUzDZjRA7fdXUtP
52PAI6xqsc4i2N0Ri3rVWRbZxdsVgjj+cmZrSaPcwE71+4bqpIryafEFbfo6RlHXdTCForySeYsU
Ut8M8ATeqIJm4zJc72iDu3NWtJv9jXBtV5PJ8UufpdmAeuNCJYzdx7Ld/IE8oa5/bIDZRGYMFZge
Yb1EUgmtU8AZtNBd/x6uJg+LsoWaB4lO1zbJyp/uelQamY4hitf043NKXRg3gLaFZ5zkcCCKecgf
8GrZZt7Tizp6SnfToAZeHvDGEP13IZkpdi9nfemuerUbKB5g13uK0vnKX5qTVj9IeVc1CDLFD8HN
lXlZBjBOGJ1tX5qq0slYMbJOchOWg3XcdFwR6xpsYmSmRsmAgL7Ea8ea9nLdnjSmLeMdWESk1kWi
NDaIJhcfyKAkpXMo0a6+YXCpshse+T24+K4S+cFv8DVkurcwGeDLUGS9r9tbkspb1eRopGe71646
jiLrd6FTaQV7ztuGC3szCZwR8BHfvZNMGBxY5XSgZCr5hAY52SUOPaQ/nkxgF4s55YvgmqzOnxQH
E1R1joJFvt7WPdoTB92f53lwlFBOvVj47oYDeajUwl2GruozZre+jIWPR5iFNmH7CxKpjQzOF50N
zEb9UFFjVI/MQHUyym56tdHg3sGxN/JZwkgbZNYFu47VmWeXhuQakC+EXULFSM23lPG9vzcMG0Qm
MqbY9cv561pcA0M4SM+ZGrrS5WQucNjNbEw7TZEyLbPdJ6cMaKjaiKegzgYFJskbil+Czw81dqNj
iS0cNGLtYCebBB+a/MYRiS9YaLCiUZCzDAXqiuiZEXA94FRVvouv/1qfHk5E1SZMWRMmuN1S0iwf
LN14kQezBpVNcvwXy6SndSFgdjCSKnRJW6vetYVVCYFMIowc6wTyRo5okxfp+elbkRWYu+kol9Ra
bJQs/V2FtfLE9DJ57G7Dvb/dwXxqjTvpeaLPCPD+CjUr5F7JXi3lpjIvPTcz8Rl/ubxDi1bqDf4P
m/jNA3NRLe4FFWqJJxhVP6bUmB8yGYGl/J5tapqohBUxCksU0QD7iqTtyeQUpiYVaxnVJxPO4Zy/
PN3fG7yKW5cxeiOFDxYTzH8mBuKrg0qOCqEKL3J1Wz+XjjFpqsW9w9TaOMhbP7331Tseqnsm035g
yv9ZdD5T+CpxW7f0AtsHtCn5KlQoduH1sjvPKmS7jKeK/KX4n9ARkvRDIXaqKE04rJYZ8LPzdm8e
vUEgDVyswwIBWu8DfYn3ONGw9sCOBGEuL/EsLDPtqaItuXcTz1PvCCORylESiCbuVda1rHsQslOg
OIz2CEGbVmKhMTR4UWiMHAWBMIrD4I4+X2vaExF8kZpahOvNWaSzjaXGpNeSoBP5PeQCuHPMMzz6
JC1EOyI8umCykt4JjJAX3ldhn54kLueNoUrdpuUbpAzypEHNipm5eg61HGKxTtFrEdH5p91ncT/T
EoeFjMHsQepR2J9y+QgYYoMtq5TN9qAwBjpcU1TEoy9hUAY7WnT50UIPGQiv3DoAi6VdouLu4CG9
UY4G5JVZbD8aLWPTydot5Mu6njP2uDf976ahS/14Pn4kOjBoQITMn8LJ5n9xq3nYbp+RpDPII6Wn
PxZB1rDBxyPdWoZeFSOG/Pi43Ips9uaGLmy2/K8kCKH6mK5RZ5CYaIZGhoBU3NtetN0TDfKgvDHn
K9Av58jePvhBR+7OKNbisAG0iBoFvgHxnlQIXkphAwAByAg3I049qfXwbZw0pVrCFi8xfdBnJbc0
KU/2ldduLpuZnFCixVCWZ5ZR+N+bw1QUgECsNT9u7G/pGiaohE5CiUMgANqQF2V5iUdq01SpCVun
OTCgGz15lKFMRUYxmGaBCpI57aYWp0Uhp0AU5bFPKpuqt9v8dlrewZLgT3dmriBUs89CJqEP01XC
hsCpmow4GCZSsEpLPiNdde+gAM8qMS/JvHqQsRV26YHRxooPHj7+X6rESXolsOc3WuHZTLTLvyjb
Tc0iuLjCNTSey/dRnXz7tiLf0CyP0ug123QXCLEed+2BMxrUSikLTu4IxcD7Am0Z37Vmj0F/6hF1
oUGli6vbE2vxyFAc2Nd3Eakv5oYmJIhZgBqAtI+MmHcfVOoZ/WU9Xq8yo08MCahI9KMlZJiEybw2
vmgWUWf9L4f7R0j0ENzwq6eFFRcMETc2yCBAMMQdIvF/eFrMiRZmNPYopWs6/9CgHN/XmWfOiZ+Z
crV9PJOI9r+mhktEbuGsb8rU/pzDEMN7Ny9xTh/32szD6R6HfjRGsK0PoXJHYfPsD1hOFjytPwWi
aSmQY2E5QglQpAUGr4/cjyzGjMNCSIRFoT6qqRWu1jvdpWxUOZ0iwsMLZm/Nxyj/SfxL/8mPAEa8
tBByk5KmisPCFF8g9Gpo/Au6YZh2KwoVfz1BWC4MNKJogmp9wh/1LHAyH7pNCsesqtytjP5jySoo
RQREdJt1UsBaAnXgndqOVoal8fmwudxB5aYREGz+xB7FbgYq8WnYIP/heUN9Jp1CLQ+0Ind/OlpG
AFpKR1v9CYOd7xUX2e/bGBfIIw/T6UIR1fVyOZcMwgeJTgCVI8n9Sd6QOOtZccLj7NKr8Sfz7YGS
FmT8etbj8tM2VjFO2qOJZ0JAOPN+0lDo1gYb29CrXEX1v7GhW9ZSqMkgSntsd2bwdaDb6HuvhAVU
9TPxvFvkDTJv9EmEO5pAfk/IiJTU79LpOzbfxEAKaVOkvNvDZFBZSO4HrPxsXknjDTbGx9njyBBN
6JacmesAy3tlbey65kFTrKH11FuQsxNTYSrBoYUDRZurWS4pUHyJWqaEn5iSHclA6Wox7ZqWEHB5
5ulvCbS5gKoB5shtDjH1jOAScZNAoJOIwpJGR8HMBUUUixzLVU50Zm+SEE+jqLCdAZby9cf5qCdz
SW2+dpw7fogIJbntqVMiWEYGKX36kwnPrfS1bTuoWyHv/VO498Co4PQRSO28bTtZd0lvh2yJj7Pg
U3ublwYfQ0/aMEgcEwYARex2bxtZlGl3c0PtScwaHBRbAaao8XShm/4StfgGXa7c8JCixHVDkchZ
HAiK33my4MXm3SGejZtmG5/R+P37XoOiAyuQkM/9KqZaSPuP9NQZqIoTePOMuer1QqW43g9lrk+E
n2WT/D2vlVWxkEHYusrtIzbyHNUYnfNyxwLhORX0+IVxn+UH28MlPKm21XcDvELl+7odLJEdwSqp
XZSx0dbnSPXeu7EGvTgU9kjE8CgbtjboJTICoGAnctr4Gps/VXZA++xOlqs8MN/e4J04I1XK16E+
ZsmwhugWTY9h9WYmv9egejQzyT1WKiey438fZKz5dUNdIVPc+htZosBXZsUD00Dp1avyhgpJuANZ
CabYPCEY82RbMKUvuk91EAKYz28M0nWb+AC1x1FHY7yaxhnDB7eNwwgvvIiGWyCQBbOQlWeVE5ux
uakK99hLeKep02LyhV/q52uOEQgeRmBmtySjdf7K/b85JPW1zR/stsSU26kV5pNxaX/gkH/yKhi/
taMIacnVr32YRPupcwqi1SA1yhmqKQJRKJfCfZApJ8nIADy5N2b8GKs1WD+1OvSOKAXBvQESPm3i
wB+DqzvA7g5R5CvW0LOHilpuaZt2WazvsYTCbqDv0zMtpYmqDEMh13qmHHMqCJEK3jz5CqRIO3d5
rjOx5bruIznRFpj19GRvRgedSwwrJtJX92wcbJYYeRh9Ek8f+Tna+ZwqrQJbQAfzmqScm4s2ih8s
GSGisFjhxt2HnEDAQB1JFJ/CRQx2yGg8ZoQIxO4kA3UW+uIxqoXK5Jh0DT00+eJLsJ7movJvKiZC
5gNmsMjGKbwYoJ0gEobReGkmG34la8MxKcLWwoFH8GiQtGm69ceJced+HNuPfpRdbNZb/BQ4rmsj
XBJMBAtTXyOWHtwl7Ie3pcJ0JbWov06MHqQcHFKBKUM2UUMwYm+S/JYjJTtqjrXUi5Bv+3DNvtEQ
JmqogaA/zc5olEIHC+Drn/nxdA1ukg8MODXk+inU3j54Jtjh4R68bi1pv221c77QRL1vbB5v0F6Z
IvBImIqKGRyQSG+al1JQY8qBQladc4FE5QkDMyN9qxE8c3GAJaAduICcIFXUT8OH9/tW5newSjrw
gBK8CYdlqqWGqFb92WTaHd+VgNYcLd3zz+Z6pvEwnSDoLCFOnWqJVbAE6G5XkagcLwob3X3CS58O
J8y5tUgz3Esyr+S+zm4nzdA0M2Sk5mtBaRmdR3MyMlQIf2SCREE9LWPJGhwIXMmcbocdut5+i1qr
g+/QS6SQNkV8J6oFl+v/NPNVMG7k/dhMSw8PhIaA/uFxgRdfores5vO+qB9PHtm0yXvtRA3TmIoK
D4oDiBhJkEbagyx/nfBy9XwD9mxYUCz4z9I/SjsK+4FGtMvFfQeSRPmSbVt2Z4LaiHGHZTUQzC8H
ok3E1AS36QhKwCImop8KicnmrNnQmtv+rz/brSUv0TNiWAsSYYRL/IzKI3IykuWiT9PZrWDg6Oau
Bgrfe8a5oMQMPA5enrhdHZmbmwXpkTLvxSqtUf8U4cX410gZhi3Y2kXfiGTN8ZnDBUDoGUPWcau+
wc8wLDvaaczdO8Eb//e4w4hx/mLTjHTre3QpF+KmIq01ynncubElePwwiEhwycvHX7r5B4E1B+Lh
XinvPtvl9NHP3aj7jpv5YFHlyd49UvozoxU6o2jy1g8h942z6MMxp3Q0A1AHh+V4rYs29yObYa+T
TvpUmakfv6/me/Jbrnh2/tNUnAeicfXyTLeLDATGQbBr+ROhVSXyWW94tv54tcUAzUPBn7qfiRqq
cLlUOM15pqXhTL8LddlEKttcMrbpg0vBeutRsNJZoBdQG0lxGNeLJT4NX2Hy6Sxu5W/YC3oFOusF
pTcjhKpooaVcAabulrt43yTiVT1s4pAfsq4RuXQ8D1Xu0TQFEXq1vcamN3ufwPXuJSCyUHmANLR+
wkrxgDmebNqiVqtZrjb+ZiuF+ZTL5Emn27672S2UTW+73Ct34EqiSizJ7Xj2YxQSNGhJJy14z/Jg
BMeJmbxoH/142EXpyOPOUx2k04Dm+QD1iDbVQJoI5dEK9T1WczjNxgz5HhqppE9++cnz9PXAsbhE
lNqAK8EHfWjXJoWY2i3UJlL2Ft/9+3ZQOanGmC9vzqTiXWrAwkDfhikSTHN/OhhuzP/aiHg5QwU8
7H8OhiasyZSrzsZ3H721FFRJ4lFBJhUkZUSG8aFC3qcBjUQfatWq/mrnDmsGgJP/NHyQLj9s5LuB
iFQZDRrre2fBvDDwK3z+KJLSvdSxWnIsxOI0P8c8kEI3l02YaCDTy1UNb3bXGPW/8+QkXi928GPC
oU1Ddsygnb34RWkUMfJL9OrzTMYmdLi74ZZ0GeYZU0/hV2vBeJ+FXz9n1Xwe7ckbf42gG8FOBm9j
1C8tEXEH/quwU31t6XEsEbxHm3fZcgzLI56nRbfpzCdAldqeDO/ZfzRWfHvjwPPFnBufqj0lTJEt
oTmZ8Wi1L5LjVt19w2UrT7KTkL6t5VIDvQEsw2eWzB2w94p/ibdpGXWH3e+NI1quT3eeTGH9w51g
+iTThKwIjJ4gY/VpdUR+y6h/98dNtEYTtutJ71m92oY2ocfavziotXxxo4C/1ANMrO8bBSv8WjNQ
kcjWn7MqoD7p1+ikg4wrWHY6jjwJU0C0Hf9dt0QuVBN86QiFdwPT4yaTJ7CJFpgpIXzxpPqUsWGL
eUzC0DbZn/OTJtbNqz2lagpbew0Btm20S7XOOafXqcMsxQ+RnAd0qU3N54xGLqpSN/LKCTUvebYV
YNhJ+NpEqRCPV0bLxvETO7Y7p76+LxrsfPrBLh36cHpPHGSNbWTdmdH3+877cdQEUKf8++Td8vbs
5Zj1TMUXNuqVdqW5neJfReRcTpSInq2p9Vag12z6Hl6055ZhmyurhMUVA32aBEnzR/RCCPuTOEsc
8yqt+/E2H90DZpUAKIis8hKvReegYSNccXrN91QZF8VwZBAHZcKqywusM44jT3bgwlI24TvTy6pH
vd3gPyKn1Z5V2ntuUTGryNOQcB0uZ/QB/Or6tRpgdT8Nzayb02bRxzDJYpaozwBVHkWGf9qVP3J6
tcPnMy9qLzUJENi1mKtk+D6iBMso4OqTZZzkP3XNI9xQhR4ZE91KD83wkYOHJ7CJxVFRdWKUa/vG
MydMfuNVVrMc4uspvxNDmLBrICZTvrSOjToSkF6yJ9mHWorA25L7yJ+I4hrByjs+ThtmUUP76H8U
asvhEdyHU5hutYJWDT7XsEc/2CqY0DfaaVo7VlAa1ZIk503TuZXmNCru8su5LfDZWs/laZCUhNlu
J9RZoA9AXXrlq81VUyt3vLZNwouv0d6RMtEEwWQA7L0xXUAvAiZMc4HlgEX7RmvKMjzxXyq4N9CG
AEZS1nSktfyCzVHWcXwxwnlGyWgaYkQ8BO4N5DiIHRYKaFA0kfW6G1N64um5k35MKh4+ijLW9379
XgCtPt4821dYNeN3eRXVOIaGhtwzoqcqMvgKI9fLgMoZt2HjYmvEh115d4Pb5F2sQs78Y7vfG8NL
OxXNE5XIUYL0JK/w71wAjb0ZMZoC/Ud5D14/hsDsGLKmQoou4nS0nvQrl42LayuAOwTMNUigq5Nt
CknWNhysJd3F9hp1W9huEHeSdjqt3ipe746gN9+eMJcQk+bNCIesVz+wS0Bare+Wp1cNLIc3NeAF
4kUDDOFIH9rpigu4z/K/GvZ5Nkqsq/Vrmzn8RU3TvVKyoPESruZQbPscQSWRtcs4u4tsfl9CIVha
6KsEl0RzjI5ZiqAFGzTVpQ46Am+oiVPu8qn1LULYaGTlfvsuaVMKZCYoafweiIfg3VOx5Yqo5SBy
oaUQMtQHMzFKEGh/ih/vniEGGvwT2Duxs0W99pP+keS6PqLbvu9HhXR1O4Hu/Ql2VEsKfXEVq/Jg
txC4QSZuDL7kqDFV070x1WOWHY5DZs7vP/YeNLdeNpQb01Q8sZpCexj7YAMFXhMRufkz9Ut/ptW+
GCWM8BTIsc5js2P8AT5YyMqV3cVgbtYjpEE8G0OBK4q6vdmjgT32jvaUn5M1Yf5CU4MEerMsd0UV
3HOvihrLMdEvclMZ/dHFXCFj424PVciLR+g2Ji29KwGIkKExOaNtZLk9VS/E9Hxwvpy3+A2L/mya
PZ3UmaXSeTssz4yc15rVqb0vDa/5b88tjYstjFbWBY+uhumaH/TMbuHIVI3vihOWJZuIIZ1DHVme
LbvV5yMfOT+pJtwANgBolydaOAK1leEMf1qqIt3NiwlNFXKWzwwrLS5iLEgPsIxR/XT9wqPs1L6/
c4zc8nmUG/s2gq4yZYPaXWC/OX8yS0orRVE+joSvT+T7Vzmf3nDVAB+1Gc8I9vb6jeimd5I5VjvS
Q5aC29ZRvSGM68Vs2pBUy7YShO03/x/vGinTU/PiDXNsgRNo4n8VZo2gSGzMi0CnR0uQyD80jalV
bazu0K0/geM=
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
xI5rRsZ8D/mWscsXgMgqvONi1IR+WUmvlhOeHpoqbkmGbmmCKddy2Qan/TbchxUow2f4O04cfAEu
JYQ5L/DafoWEAHShGyHztGxj4EyJX7x8yqtcAWwgcJlMfy/2Z+sYHVx4ASnUNZeQ8HXpWibYIZuP
FjkTNuAr1SrdQnqwhH5cviaA/5OheQSigRQCP8RRQlRyBxc+biSsCZMpGISZFX2CZjSyU+7V2yWW
ay7r6zDWmMmDZjudTCI4MmCNXIWpp/bhBBuYrBSF+L/5EsYX/jb3bbE7tKSBxKDVS/NsrCqqNgPq
LE6lSb2eW+8BDcfgsBxnkhOXEUv0U/y1UADlGQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
kt+7rNkOSYrcXqbgq36Tjy1mVNbqyEaJJcQomY0hj5jTsV2loT+ykCqTokaSF04RFimKeTBrbOMs
fGmY0J0Y3FLdb9mRm02LfOxlSlD1IAUzPqmK1XSR8d/4MtempkKY0sPLjad2NV3YwFQOuIgbOEwQ
WJexgoWi794m/yDoUFziRVt8L8gAHObe8TsXdCCkIFw1w5BV4qiVphOfsBcAFfGjk1h0eqKL4hHd
+knMywKT44w7gE4DaneMKpcCfQ4X0hNR6jP67PdO/EqqXFjgnAn0wypmmiFT+lBYDb/eP0n/hSzE
W8aox1YjaQtyA9zwXG2XZMpfhHFKcSJlD/u2/Q==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=153616)
`pragma protect data_block
RvX6YNnGq/QfZrX3+SpkwDzMRMPNyB83XtyOs+h+gSiynn1XhUeSuYChhjzO2tVQ1rH3F/vCPrla
hD6VUALEq148nibJmMdYwv3hTk+sBmRcjCK49iKFYZ/tdhMSsIm1BIZrY8EQWICi7teBeErv3NJb
dWXAjbrToZfLhLs8dbOHQ5IeERmI2jxMHlIDLlxjLEHqV9ybINIEoYCUNFIKX8yrNAOSiB62AVk9
F65vgb+GThPHJp1sNpOWimfOv+/6Oo/W6BOOxzOHMKJY1us6t162gsKUU0fWBNrCj+vssOQq7SrB
crH9zn+iMCxEK0YZzuJkmCMWqZ7AZwtfRM+qEZNUA00xy4hADuAOa/xj7enRywhQzcafss6zoYIt
1lhyGaSALH9yhQlAkHYu1D0CdjsF2iZjIP5bXsPkxW9PLppuaiXqPlKiBsWHlmqTgUB8FnhBe7mM
kFq1zezqUIAflT+m33WmUalXKUHOqtdd0635eqO5k5eHI0wiUneaFAdCPFejIHyNFPCTvUsYCHSX
283+wbe1rbMZ+2ed6HIEA+kaaIKAxO0MLoXJGZKiTILw/G39+wS8OT5Xp5tAk5o2LnWbCSE+bBS2
gJ+5EK2PMHiPWhrKT6aXZzTlM7gHQn2cd7Jclduq5q3iY0AL5/AuDwITwSYQH0twu9KT9ez8D6tY
OTgXHwVBQVIcjZSk0pDezZfH41cqEAfu46BpbIxWq3h56AqwZ8x3EgOHLpvpSxxklNmRWyP2EywL
hh6m5Sfl84TE2Tr/AszoeaNR7okijFln5rsOGxKv+24JvMmMM0FSuhl2aSQBSIJPANY92jF+/+8b
d9vF8of5V+KIeaU7PAGqfuxhBlqWBQ4zcc1OvV3kUs3LxT1uBKtT3swa3Xja3JwFUolzJE/zx8cR
z7XR5sT319n6K4xUvhD2naLGMsQ5G4hHNsfQp2+wcSNfTtMsTxqiFGOaH+BX37mM5gnvUr51P0yb
yc/SNgXBvuBEoSNyNyGjUIFjxoLXekSooos7+DdzGJ8n/4NBrK693UFRjkeGOx3JDi5QqThVH8Kh
mJ3tELLl6f3MBhJcaaBUo9AHuCJyTtyLiS+i591GJajt24K1tilzt1/1PoF81irDg54UhB+6aJCG
fO4wGlJXfPVoFFbzGTjI4OU4gKQs0iLD7wQZ3GztTYB+E5MqY/ghXYQ3+u1AOPqv8e6cuGJI7m22
Qc+heGoOMGV1AIgCZFnNAOdnEXSoeS/QxnKGDaA8btg9SltrG/kVfInMjJkd3UvFpybzM8j9zs4i
gLSkVtdoByly+OKTzHRRPrDSoMtAVJ0JmXVgqkVqJjfy6DfDj5HrwLQQx9h5Kdfam4Va8FNYeMij
spsIKGWJ6RcKHZ40nDA+EXXhyD11fTbRhtOc0ui4+7EjzPQhuU/cMKeMSm7e+OFJ8LImQw+/Ufq8
qJL2dqTLUpgM7/BGpPcVIzj75dPF+fA9CELZ8hPE5l8i1ODEWil+6/rgkf7qIzUVCHt43ftXHjD1
F3Yns4n7pkm+hJ5xnBas7RRxixizD9P3kSWO5gTMuvlm4M/VjAtKqiQZQYjkFkTg+FG7I5rlSaIV
4Vj8GyaMp5l9TFTY1Bhl+pyN5PVzhqPDCh3Wd+SGQdgoGy9UKVGKnpGpt5978QaO6osIJpaAZ1Y9
h1qeOJ0WdB0RRjEEzTGaG1Wt1r9Rbzq3v9hMR4ILVkNqw4q+6krIiwTFgZvzRGjDf38b20MTirr3
R+dmuIMn9lgkadbWSBfV4mgsAUTCdbENmy1X1EMJLx9EqhCQkuCmCvZ89lAwfaDTIDmIc6oX/4Nl
UMAntgNyIF0s0IbrVO8xTbl4fSUohEGvrjpiUwcjgj1089urUr7Y0sCmZslzqBHwnKj8UQHp1PvQ
0D4AeMvJuSPOLCcI9r3UnwChSJ+JiiwfHwZLrlH1/hWe83+elsvPMuQp6Usw4HuRkAgKV+X2Peo/
p0N3EQaYbeTKu6usXYwNjwYFVExOeEFEglkhmFT39ArB4zweh3IhzbVfH5hVG57JUv1IlVHgqJ1i
GILU6iNao8AJRzB3Rdjh0MzFVsRaIPGwZ/P+pJMAaLFnxYVthpP9RgEl3/zIdDsyl5v1iWta6brM
sciKYIDuLPBH/hEI3RFwjFSZBV+5vW3PgPDY9DBZjH/FkWm0FDxWfsgUiaUdEMB/mk5113EjRgua
dD+8erOdgkK5E0zKrSO3c2qW9THrbhqL9LDQLLwzki8sWQY8IBvqvfU5ZK3VuJatFwFJamv50lEg
A/5tOM4vLCVq7Uioy1VjGNVG74uyMDU6vplCtNvj6r/9tLliEoD03dpoyeGp4URJoP+D38c/k3Lf
TgquqC/Vv4+3uugECDUb2oqUN3WoG8YEFq2q8xRIpXaSnzFapG8ygKqK/Lzdq16GOi8aJ+AXxlZ0
yHtHBBVt0t26tfGB3tz81kFRL5r1lpIEDsa37FHzOU0x+TMoZE+9EfEaQ74IYmcB22cF/AxD2ACV
W5LqvppKhDWzBDfOAjIY9vi/p+3rNRdq8BnfuP+33O2bQ1ZOa9FMmfoV95DmsnzjNyXrAvmdLBMe
DjZTBuW+ZWPZdqbug7zqveCmyamASgjP/uEiPmiUjHvyU+JYh5rXqwHDYglUNfalNetTq7uIIDF9
dTMW31JA/nwGhRKIUlyObCSkZA5Hbtt6JxHnWzlMicupJgDjhJcYkGrXBzp/q9UuUtipD0hcmpRq
IGFoiZzjL9jcDlo4uBx++6izB/9RSoyBXsNwbbBKARNePk5Z36DFNhXfu+LkL4ebnIHpnDUVg0Ds
klgivCH47cttZZZuLdz34gSwO0ThdhmWEosjfsvxE6VjHB2zWs6+Zdeec5Ghv9j6uQq4Jil5iDG6
VFdPBVWk86d/OtQSK3t8U0lfEWF2xXsHHb1tR/dy0RQ8kJSJhWA5VVf6FIrYtYxx48Ds008mVJoK
N/R4emPdyNuWxfAcO10ork/Wz7JQX8EIDVpz2buGQhHsMnKHGVvsswEVj94wRXLBEzqO+r0qhVJ6
PsEi/dUKjR3j80k1cQDliJx3d6fpQlK7DhkfGnjqumwpa5aCJiprB0F4aJ654lYFVXpvtQe9pwPK
MjBCHeSGF8QJ5MQT4Xg0zyQHuff5CWJLHrES4qWYINNIX0QumMK4epiAvUj/d4pG0g+Hkcx0qTxg
7k8fXd0KXF7k/Nu1NKskDGGLhXNPrP3UwpOmMuRMMF67LtXJkBpG/QQmoPFaKIqGMMuhGgL64k5I
gtYDlhI5OLXNuDYBy3wjd6CqhFO124cBC0Ph+jeH2H6YnCJZ+9MEqlHmTc96Oyrf60XJHMk3UG2A
KQ0Trtgbp6V8VA2hPjfx08lX6/msAX1VzNpQaJzKZsfEp+Cy64atT2K3+66BVCj1aCdLfQonCeJQ
XpAfKhLwB36ErQm4uPhaSoCrrhaB7rzmYVt2JJxexUDtNF7ilj1Xt/pXnUj15AEs9tcB6u2ZLtwm
lWS8t0wUNV+EQjiJMUk0hm+tDT+8DafWG1IfF5Yctjb1WobvgjJWyeSyaO5PNWDayRbWiUcW4Cry
4X28SF0SOnrv2Bh1fNIKUtS4Iijvo7nI/uiRCFdaXMMmoyth9RA8FU+o64VxERqfr9beL/AitdjA
Rvonur6rIW93o60tmRAc/7Tn9ig6dCN3cIP4a0NwjAUDNl0Bs7A1sjHEjU80T7sB4CtHWbEmYE0+
pi6yCg33GXkbJp4x4qAO36ccefEaXrRm6hDvKLTrQtG2VYPbds9F8hKgErDId676A+xycLuWqAKy
mMsycEpOWZbKseucgKl+z9XceqSi/vVMiIBs1XNRXrvnieeLkpWrg1ZTR/1ml1gP7k9hUSSZyT84
xd/g8M8bL9Ux9XO6DauO7wg2G9N/+EoROoJ6jfrs+FS2GHuvdn54XQpa5v6dSkpXjwskHiQ3plNF
j8vdUGL47abfkjcul8Ww88LpxI21W9bKW2fJfgSNBa+ROmyd+d+guGlymkQzs1kU+auTfyd0L3oy
EQ7afX6PB/1PO1jisVNKiAr87X/EUyg5xH3NvAIoOI9NRg+ImJQB4LetSi/5E5wfUGbJ5HzqOyO0
4SrN9PLd8pi/7ovzNOJRn3Up3Xae+2lL29ubDb1A01cAWvICS0W0+RI9KpxT8fD1BuWVbJbVQIVX
iJOpbhLC3atSqIgqUK7RHageZh6LCw4kXPtBMn1GhPradI4nf2V/z2IflC6c2vt3QUWoi9EsVIbN
Uh56O55AI20yuqpiaOtDPjxCqF1zcM7iBRfSXLcDUOjCduJXlPS9IMT1Zo9mDX4PItVNEmhsHvbA
cTxLjuczyfcWTsDDrdR2a8iu7FdPmNk7Ozf+B0saXzUApCcohlSOsaMGJvo+96uaegxtc8IFSSrS
ae0/oZyDitOmTEl82y8TBJPMPxJKAeIVvWtFg3z/eJiIFNRJrc13+u3WPYPUpllnDdLka9H5lRlc
OFNZDcXEPLPCn0HvT9BVFuVP1ZBonesHLnILMDP9+A5MJCOGZ6BQ2JU1dFoOjC6eZKjlgiRADH9y
6H7EFWt/++Xy2DeMYcjoFCdr3S9BlD7zVbjd4NAX9HWFfhBWfp4v6ZP0Fbu9YAY2o8KM6NNtXBBo
Tp86QVXb/xL7gUn5xI+FG02uCZHSLm7pgJhbab+tA8ohHdZys1GI5kaQN2OVeKXGUsI7HmyGNE0a
ogc0sZvsXSchHuq7BZWRaDk7tbeNFKSURCRz2Y6Z46YXVuA2+cOC1oRaAeFGBR8/6l3OViXkD6hv
0DXpBW5SCKdPb1UFEz1LU831KR+CU/sNvG+fa4sMig5Mq3piuy0upqvvX1kbqxoEajch4Me8aHsE
0MctaUAlO+SY5/7CHG2eWzii+AuqtDGrRhcfvL2/3qqLct0/Wxk2FNenNIJuUW6JKOHQyMi74r5L
IT/D/Kg9phVRtIbLgV6AzZfRCS+g3gL8gM+UXn0a5pxrxZTEXnopsjKg/CkI59AMhTbyElVcKJi7
51VOYWFc8NIiSN/lJlJam6LBWSZf/mdPRE5XmhU73EfRK5XH7CkVbTM++a/Sy0lTEpCUEvIPeCoh
YfIGD3TYV9tBXfbYuZmWSh3HGiC6i7N2gCQQMB7f3euB021ZeRZB4yY/t4u/1jOR1D5U3kNeBCtW
TvT0NYegdOjtVJFb6Q3a6bm78AffzUtBDOIKkuWKXivJxFufImYE0Y1s5f0dgaLNYaLKb9OMT99t
Av6pUSiczKtJQAyGt9MdKEhujUmAWQD4AIDj1Cbh/PfqHpgOb8uOZ8xQbnpwbWCVUDZ6/8zX9eMt
BuGpzzc5NjqzDVCsn2a+7jVyD8oZlhAciCsa0JnKr14NGtW19XJnNT5woLyWWJ7pCJ7kC8dw8lIi
s4xY14e4HCpXhsDPCN0F+kSI8YDg2/A1Il7NZlPngxoXU0DSi+znAMRY1QGxvEfnBlr5eWSN3hK6
7jMxH9PBySQtwrrtmZHKThVrY2uQt506Z6joT0OMj5Ajg1hUKrMhWX/vT/1Ovxcf6QFoSJoFyQyJ
Ed2alEN0sZAr5gJGRaYRtKumkGr/YKANELFsiucHgZgbZyidCQzAJLRiGupNa7v4Mo3BOuSUU2kh
fwcm3NGivN/akF6AFPx48ls74bAq6+n+oQnZ1SIs6b6JUCaXbAwcmNZ7rQS2W/7HvqVBY2Ch0QyH
xQPlclLtBDnj7SQL6LVPyYhokDZnGl/wNWYG9AuXglLHAyOH5oJnjp3kUnIYY6YGgaVMzxoN97KY
1lPVPAmk9ZSuHgVxmdYKLBB1FodADvMJEsggXckZ6VfBBRIgCSbJvS86mMQivWkRMdvvSJ4yBJcO
ePZin0Qp50KGKOAD9Ms48HoZgWH0QmabTMQ4LxWgrGCpPrxhJcPPh6YmI0N0E+KKao/ekqBT7sox
SDFwJBsTt5Fc5t+7PXYwT7lX8GT5bsBqnFiAx6SZkdFRCFM8TClJ2WBCJRY86OMIcw5QQvHNdGsd
Fq0Mn30jvFbvi+0+IOKqfqqmEKlUuTvlU+u5JzBYj1JrM7C1Qhw5KdXwZBHEsh7PBPBaVgSHt7tK
PC7PPu5hVbR23SF0DT0A6rovMXgno/F/4mnugbnrvT1OUKtbnhNdvUzIJB8b00Ii3qRVYCAWO0en
09LBUE87UIJ2sVwSbvWEE+bTK1HBtyTv0w6Jy6I65tj05gDDqt1i4URy+gLtVBTEF6M6m4St1Ra/
Aie0D0VZE5nf4OCOX49RuH74bGv8kJtmmR1OXY75UEWiord+cksN+/Wfe919opPuYaTMiBsuj0DQ
hPwftZXT0Lwt/lVrycwiR8I7tmlP2f/u6VR5rQBONt64fuGdlJTHQ5uO+vkkdYTObBr/FSpAJSiM
43VvJ4piWLWu/BWmgqjWLeD0tyFj58j3thnnVEsVOyhIBn+2BZfjG5g5ryeTWCKlTfCyuZfWdf/H
WosR4KvjKWya8NQcrz0nvaXpjDAVOakGP+F4vXg6U///1IcYzZDJJti7qDDWZd8lmnIJFtB8JHL2
KzI7E+t32PjzVEs+CdTsMcYboA98mRccjOlkg7utTAuRnZcFy9/yuH4qW/ZklY0RSR05Wz89h68r
Whfr5ucFA5vyvbcDgIf0KbMUIyChoHI3RrnUyoalXwEq3+AWj0+ISzbipFVZq38/SNYKiwH2GgKU
8Onn0EAf4lW9EiywPMfqpQAFHNYZXHZNeinQ5ELV5qm338Q2eC5RBPhZHuyQsSyREpTc3Imbd5AD
xEIYOtpN85BHdmXX+eJfIznqejeUphxviOG2JP6imZbgJK/V1ln45lQqNIUDJi2w3qUyqsT5UCev
JKNkVOysMBnyfy9EeTPDmo+OQNSdkjtTRMSjoCFH0UIDMsB+w/l7zYpDzNO/mtvqMAXZOw/5V6fR
KaFwbl6qBFOI/PuiMr34tAJDEYDXbO8331qEmCkbi1yimUmM3H3UQikWos3qfInflUVM7Ma7AdT+
0JaQLxtK82yeWTSGD8V4C+U+g2CE33gf6ZMriUeWmFylRtxhpHSNDucKCsBRkM25hEm7+G1MdKZA
3Zbo1wGcKTesgRJ/bxdJPTQzbi7o6jXlfzqWYJ85eYpYY7VOioseuCzeulbj0dsgp5IIrJnm/fHC
ZF9nqsgW0Z2fdm/dzOLetwl6iD7VONOjmKQBHYeTzmT2CL9T53rO0vAGF6KgcyGp6PzfRQWTvPhL
7YTfCIJgw+07JsVRvKXPmmhRHDLnIR6BK2WOy+ty1lftAX0T94ECFfUVJ68C/LrKCxztHV00umhj
iDNYJ2WoVyHdFt7HavTU2iZuqEimOcRCyeqrInPwwbw1/13xHAoC1YDxYkhE+IIZ/fzhQhjt1w7V
Kwee9GYyW93MlYNHJPkptJO3k0ubWDbfDZ9SQMwdOyb9RZ52p5m1Tnw+O5r7T1oL4BPMevEkCqPw
tczbZdYSePWIKbjWb5nJBTXJq6XPgnBIcW1ZcHkdnerzllmjoQelGNrv4a3nBAjk7xqTIC6tm5O2
91lJUVh9L0YAohcZmxXqwahlIK7mDDFPbf6T2d40E6w26SaTJ9hFhjYB5iGOrgvszBO+GuW+YQ9c
kDeT15yjrCgifurCi8hezGLI5s06Y1IMy4UDZrVHd4UQ4iWfftItR+KGGpv933RqB7O1TyYVA/aA
vBrTztlIZZUX18e8mjoBk3pTRfpy8/vhULEfZK9TMxD2oWxTJsvnmTgkyxmRnMDtLL8nFauYTLb8
+R09a/FNLtg1yShwvI4GR74YR2DXDOiX5ApaQ7wBr28ZQcU9jshDMWlRjF6YrMFwVHLJe1E0uKbf
gogIgOWkgGcvAWu7Qq/A7ZN4y2Uu4i/wIKms7S2d8WjnEqxtWkJmBj+aGYhdtt8pEhvjVCLhKslr
Vu2u/kuEeaBBYFcdzhjqc+JkDYAZD/gethEMkqgEd5sSp/PNXEA4vBzgw20GQqX09sjmUyH0dhku
Lpo94JJvQg1aNeTj4BBDNW9r20lwolWpVEBD+7U+jtMxIIH+wZOt+u831YJkAYLes8ebQUmEKF/7
XOjrr1fAMPHnyh9R4XdWWSvtebBl3AWf1c7Ay/BA3SAX4C5BGLpIKenS6kkKCuNFijiIu62CMYvd
b3OQZF43UVQVzgD+61ZwpOemf7a1wAznTViFQTvvZ4C13W2f2s3jwQos1juxHIl4LuxMepeXHHVt
HNlBlatidl9+S45fMKPJFmyS8tp3XDS/FwFkoJsUqKdvCRMrixK5sXYi0Djn/svyLUikREJSxy29
hfW4HpSwX/UECVuiSffVYG7Yy5tqqn9Qi+BIuImrfo0KdniS/1eSj1NqHFeDSVC8JYXh4+yUlAYE
0BidfXtomyg33KwPOVHo5TEXa7R+8Ynof3GksuJO3Xm5IurCem3IThfo9FO29wrIkZPprMr9hEP2
VIb1Vx0pXz2DenA6kNw280V663Ew3/ZIdUZISPW4fN1b7XUd+EVVUOQpw6Opu9UwoZSyk3413XEf
U1uqnPvAQ0CYC1tMPrw+Lj+kdKc/fwX0yIqfPtHoA1MmpM3KhSMQ18O2VJA1qjhpvM2CWgs74eB/
k9h2bmGbq0JHCLcTwVP2pHpXAuCq7tQ0kgNsGSTlPSJqGa2ngVn8VNcYEwdujUJA2gM4da7NV62+
lQeii5RJHC0t1jk8JpX+UfWzUnPCqlnb4U5tR92zZOSyNUmpVmT94JFCe5Pkz4WGrn3Coz8I/MsX
lk/AlsZH0qZzh9a7gZZaylHBFx8LQs73toM5WKx6i1UrF1g27LbvdP34YLQOQMtOvgqUIcJOz7Fk
xVKZWRB2+aIpERX2ItQpNF3PSD3x47/KQnvL9KWq5Y8sWOW1oQG4O/iny07woGv/K7LjpWXM2V34
Bkgqo6Cbvl4HnnV8Lr/PcDtsvdQZWRWxEaa3fxYc65LpS8yAQ6TY5K41cCDjDuzo4UMFsh9XoriA
vqgVC736Uj7yn2HONRKYpHl6uBpmAEjRkmiocPKAIb/qngPnm3fWvF2lEcW76P1uDim0w8GPFkmM
ALh5KP43iPgHFk+sSZGit766+i8ylE5To1UJGudcxyCwXXV62qv+WCPsMQe3NQqJy/kARKFvkY9o
sglkl9x2V9WXpAzqGfHDgDOJ/ShyVIxtLaFVWUsQybYEJ+cmdlHM1ZS5WXj35/IvgW0763XkK+Qs
6hWK3dQh2bVxglkuv6ZZ94mER7TZ6WOYZpxpW2NaiGouSyxJYY1M/+npokkrsGNtqFkKAbeUvX/E
pYscjZKedblRoumQSCKnu6aWhCcWHAfRqFJ8I7aOdXhifp44XBT+J55HD/hzb6SXvul3IFa4y4nK
tcXqD8kscjKRhi/7VxNF+wlIdPaurCfS6eUZB4Jg9vDDM9zz+jA4BKTshBAKpKs7W/d+OGjZNCRK
SDk6cbw3yTyXY48Vx+8TUpJahLR4oad0rCTtxfkQruQuoGCSnLQKtnwwqRhEVsKHLUtOwk8nNIAZ
CsbCHRFJqCffqAHoP+xR8KrrGo8Pqe9YJko5L7VjaDFDGKD4cGXFHTsEIQAn2Fa+Cng2AlgHJcNr
9IYY3L3K4SaAvKC0DI7cpVBNb7LJevu2oWCUrOuYBlP3AjF3kV3ADDfV3u2c9ubckCbatQF3hFPC
cJ8kC5w+tdL8AB1ne+qquTgkEW4dWqIyFx+/rZ8BPaHR/z4ieusfnPWqGaXXU8Ae30ZLIOhzGypM
9uYXw11MRWVA9x7Ian9V1HblaHEHA1dLOiMPehxQYyKmczsGf14VpCfuIdxdSBvduKxKaDvwfW0O
gksVPSJO8UTvvLnCIm09olpDbggR7v0Npf9tunzLz2HHuH3JkoZDCfFHkhyDhgoEpErtRUFKicb9
WJmoyXbI/d7KkJO6wwP3Q2tHAZgMova6a8+sFHfVPeKk1w0+jtnr+RmWCJUDxEdIanH1vmHHWbV2
d3k6/xJzzNbs20uc2AqWmjH87jLgsbBD+kXqQyoVk5cfoH/SwTsp9BwfObaPnJYrOTltX5o6Mtpf
a2CfF3Z4CtpC1PIOiRRQqSQLk6mGEFR/xCR1Q45fgIx6yyFNtyrocV3TMA7b1dGvMpVAJvFr9DDk
TYRoStw3XAXYtHu2C6Y2SjGY/CyZ6Jsx7rAwEDRpkb3U0Gsj2IiE/y9HAfg29HlJZKJNqxLtw/AD
Th132aVNIKri2ilEllisJjSrF+r6G1BlEAwKFjiEx/E5/TMz1aXjCRDU0PEYYt1KVvEJLlfcarhO
L1BAnCZCQ9rLwO14X+6sHhotJgPS5BhOuRu0u7IBQaOI1lzKdy/PFJ0e1OHPe2+welCXtSiCXCER
Srecf+XgPdtS2bj7CLkuilpmHVlUkDv0IRoQFP8vtf4WHfjX2edxIoitMcYKv41qyOwn4IOtM+tI
sopLXl15wupBi/aFoDuyXVizhX5vTiJSrI8ilbnwpCS9B6cWtfNRnsw+OvHqBGagQkqN7ByAa21o
suoLADeTlfxkCePEKmC3rQQ3Xw1TMneY0vNcnXPSPhqrU2c9SUgxIHp5z8JnWCqIh1DMvybxZ+Cu
JP/IAZ73ad6WUWylUr3qrjpUJfbPFuPTQHQUeBRxLOBKOSuTOM9sxsn3rq+0ZFbSaa+RqPeOcl5C
9EKVmreDrstJx9nS2lCJ06BZdxw1V1ywe6Pwf15nIbqeKiVCVLG6KW2V0lVaHfE9sP7DFJhrOWNN
72JdQ2MUCDKABqpTLHWePhpZwY4cSso58+rpAnBf4rtDJj5XwX/HO6/LuBI7GdHy7yrETgpdZC8L
RASqKqvqnTAVyJUPfvIFfW+1OtRes91bIkbTckX2mJNwk88KS4tszgo2xES/M0BDml7txQd1eZo3
owNuR33Yr1x61rdgbs/LgNYDjnCc1vpBxf08xKxr6rtkQI4HSm/VhfCuBuBB6NZbS6MiYjYo/4yf
kHP13COYV8nOgeuF62Wgv40p7aZ6I8Yu2ntvb1sisWXBu1MAr19dPZH6Sr6sZO4qg11t64fzLme5
IxHfNGcc4M6+rKIj92YaJ9rxlUmnOvCo7gl+8rTpTZ4nnV+NDrGwWMw2dGW7myKLO9LeGBgPFEP4
mmPX2oW069QUJOt2GVah0NZuLXwCdfOPMlHOepHL34qktff1EqARnDIKYEchyP+J1Iqftj7DEx8b
o/XCR6I6ndbl/W2hLo0oP0nGfja1nQJoU6Q8l36zkcpm2Wfud8Cbf02gtlY+HsW+ywa7XRH3Dzt/
kVTMqZqU69dSok15FQVofQfHAgXwrztQVwCi5HJCkF4jXAf0oLdSQNV7/pmJBpINiNx4+FPJydqA
xskX+GhSn2h9X8uP3zvCsOZVr/AxMniby2JMpaHrQFZszsmmxZwTmdZuJt8wCvyZCqniP5STjCmK
JMetDZ032bTt5QF+XS6QKEfA/sz1GqmPUqwi4uYK8PPwD+vLgaQ067ZayFksKtdSHXTsOQuvf3d6
tc8eiDgAPV9GqdkXVP/xF1AndzrTMqeUZgpiEMBe7gxIRAYvV462i5dyyc9gNkE05BOY+JnpwaFV
fGQusPloFzC40yHGuA6cldR5llqzVHhYknpCPVPx7KSmUOuiyMhXukvM7fmPI6nKFV4QDx5BOWR2
+qt6MmaN4yTzY7nlz7rB+Zhc60iI8OCLHKUYYL2VXNt7gC/FlwldHxVlXpF+geDeUXHH1RsuNsir
uUgUZWrr7pFRxDFaBH4IqqGOVlNN5mIZ69eF1dI73OPwQSvvtDJrliJ8xjZvncpZ9lznBjg1ost1
g810W0l/onDAjReKQIQt6tIgK0lgKxBe+Bm37wrxBu731bSe1Q5TYIGQDMOtqYPLByitcRDCZgAg
iMa9dP4cXw84+4Jgj9wW/ayexo0cM8jX+W5bjnursNxYUtChHk9BhjTkSi7If+qLJkcUuHcNcNKU
bR+qBikxBQiTgDmTcj0sVWsMR7IGCL5dzZMM6Be6C2UAVzaE8prtAjhLjFSKDlOnXdA0ZViea1ly
iG6Uxn/2NpR5CFwUlEGVz/w5N1RML5AxDOFLpoJNdmAQfJ9DnTJbmL+T1nJzmxUPRuUtwijASABI
GzQTBHvZQItoGUJnzmwduGMiQdYPg1DMKY8bmW9b4xGjF9wC2/Qgo7VZIOgvsbt0KpeIS5cH/LaC
H4CEi2zcH6Ctx9gyGhcU155eZ+1y9ugUQyuCKa7lNh292QaM07IWOeuEm1lFMOLpjQ/ry7Tfy2FD
PokZKyGf4PhZ184wJGCtSlWPg7XRLwoWxiz78W9Q6KzOLneZzl9nsdi7HzWo+g0is5o7wRO/raII
YSAC8yi98FVzSKeQ4xfTPHvOVAxV6BMaTs11OR/0rMI2fC4OSCLP852CJleFbCS6rjnI0mBLVXJ7
/b71kXCBAJ5xKyzhRRkBHVy//FNHIXy5Q09bxJmwJG7cAfVWOtVZlYZm0g4eKxCpf2M2aXiwy4rW
+r3Daq14eHSJKK5k2t0J+xVyU/MdDfEM3R8qF+h63OitTZrWUwPWVGfztoquYNUt/kloqpT4B5v2
kd6NfN279XQaESX5y4LP+l8VHjol+6JJvPMb9HtWeBDUP2R5AkmJDnjZXAyvIQbw2Jqh7XGYsQ8g
iCGtfyS7ut+useoSXR9qm53QRvZRVC2F4TilEBOpR3YpBd5iQIcWhkFYauTlwqCcAMSVZ0QJrQI+
lKnvMQSxfIZrqs0ovbsh74ZElqN9sbK8I62l90sLS6R1rKrbXZX4pW2ZyXeLAmue+S/JcqMqJZ5N
tvCqICdq5rR9sKdhf3YzWDGo6zt6sxDggVVzD88F7dURSUS/+pHaDAa3S9clNwG6Pd0IjDhjl175
sEoBJRyVugbeRd+7NDBqrhWGtix9M6K11MzeO2HupmKs1U1peN6maPGJH9cM5U++k1VEyB2LvZKN
QJRopH+/1kYOagj5YS4cwq1AjXQoACzQKivv19z3qN/j58E1Uzy4Bn2Yko6UABsoklO9vDRq3pWz
FbFbvqz2qi7J1XRdL3vEFDWNfkzt6u7WDQUpozumAM0ipJhlLSb2LIhF8CQb/RjzZvGP36o2EV+G
oDCCFlR4Hvae1NcppupBiA9xFvl0alqrJDNN6uM5lHV8eHVa03mqc4t2xgrNj+wUebvv0EYZmJbs
fQ6F/s/y/7ijC8FwsQhy3/oEfezY2I8cq/ghIQPW0sSgvULCVQ0UDrBKDWhsu7kqAWzF29l41E+r
/FeCb8XiZqyw/SnSlhbTEumCSbtXlZYc5CNq/qGEu1Ikg6/km+tnn02DcRTO3uWV5Z9BMpmQsLCs
2hYYl3mcoM0StLwJ+RFBLEiUg4kg8LtPQTPyfv94pIEF9MLJnQh9LtmDXNBTE+ZZNuSXslvKz7tt
xuUj3VisitW99rVsv3R/DRzkaJH2KwMuZlx+aE6hkgvLhqdXKpVQEZmhj5evzn6dDk02syFT77iX
twW5ZBmptbkuxS+ku3AhhBdSWalRhf3sCT1zx+G0e2eT6Zvc06ywZc4f0oZs6UMKGGkJL2R1jBHu
Qb0Gz69IJpDuyQI+GvLcMYta+iS/jUHLEtdYa5P0/doVOWeMVGtsjFPxXYTMyPwtPgnxhC0fZRuD
IrmZepdmmYLfR6scF9GczKNHSYUxoXz/GGtcqmun08N7zTllsg7ACyvukMERxy7L6xXVcbjvasgM
xetHPr0kyLeo8WcssFhowv+BVsb6zhOaYGVfOGwyeNRMIoRS8GDJfC4vdLdPknfQLEvAv815KVpV
McIm1dienZqoXym6/dUmKh9jGz69fDzOpgMjDAnzsPQHRwtczrfmVi9Fvok/PAiOKJRioKUyMe8+
lwpc4kGFgczP8pkewCHvIm0D6sLkO9a+FmjNw6mEeymQ3hV5qUz0sQNcJYPJkCXiXgbMGMZ5Xml2
yqGm0WbXvZufAl6lNKit7iaCdr3DVHaMFGRuDV2ulJeGR/pzO6quTdA0FsW0Y6JeAuDg6HPSBPNS
9od1vUAHlw1J9luH1ZDeQgJudNtu6mr72DgxAifXVM6cd9mOuJRQXBIKU8qiOZdXQDdgLGSiPnM5
tknTZHt/JjglFBYZBrxF1B7OpHKg4Tn5Z3ll+60nSE74NYfgjZZkDd2aRevPJTwfarNihhKuALdb
v+AKm/nY3Z4YIK2VLJGkeWxw6trx6mSjnqMaBhiqNHLHKg4Qc9kLDb7uJvJCN8vR4RddIzyrXWZF
xanYWG3no3GTjtoDNEeoiORNU3NgW+7tQo4U+YNXAOW4NW+f96UM5ky8BOUsMEn3it1sYGVe4etV
wdCYswRPen0WieA0Dgj4LCoF9nl/OH7r8JNWryDam/gXyEdLsUKVka1BrEESw3THuMKthP+Z+OcV
93Ql3RJswm6McEsHSSxwcuWB1lrZ2Rwfgwgkt4OEdnbFTApA7E3/gl8OPBChqeC23dfuH5aM2W7c
8szCMsgf/SwVkXoHgHtjZZ9ArxG6vgscVEbfK4LRS1dyt7HjXY9RSFMJY/fnzlFwxYZDt62YVZyS
WHrQEGU1GjXO2aM1rDin+3g2PyrfOwD3cwMGfaD3lmTsaSxIaFuO221W+CuigAasZ4SPJg7gz77+
rzFPKAIUePac2A58fYWuT1OrOZ6dG2wwpbhqgtgEh48cTgUA3uxLlbR6RvGgreiixTyx6XrUJQQS
NhZVj/4ouWr7fib9X6Uk9eJ8bbOoXTYqBpsHljSLdb/5053te8pN/wlgYSfH4unPfuXtA+c9Gdwt
os1Dr0DfZ6sCeuec1y7yU/TMwQtVns0Z1Y3OreWQHv8fGBn3xxJtqMN4EmIer5dJFygPCNNjX2ll
fwRjNYjMLXRJkVLdoKun4mZqbWUJIj8CBtvnIyOArjBfwqoKhMZlutAdXtcbDZG1fQHD+7/t+iBi
LFWpY+RmOdwbaDTnMcY52J4q9E8XDaf4DNOZ+C0FDMw8SlyY8ScInNJwO4rOd6HZ6lmbqLRZNuC8
qziUkjNv1Z/AzVO36TpzEDO4Z95OiyxGFQ5NqynX4lmqtL/UaYaFADIjKA9I0sEIE0CijAWnPNDR
kmNwXWY6ijGt7etycLI+7JxHNWNKNMYAl9T2mFM6zSKFebyZdQ5ixIgxghrfDim9rbmlNrsaKwnG
dGVrTy8S9PcN4oVO+dOkZQQaroW2HN52E98cHBrQQAb+FjEO3vq/ZvwOF+/AcV003+w+48bqR+Oj
ZFA0Geaju1BvyPWXycuFE0HxBNOiDnWjKm25wrUdMAsbjIO25ACELRMgN1ezrnKWwhqWqfXyRSeZ
1Jonqjb92CSiNbYH3TVHhtmhhxp6EimbvuleMCrLS07mXYdD9tZGuecfTy1PB7B2eC3js33Vl15l
yAprUzWwj1M3qLGwAlgWSQwt+acHdCL9Jp9zrd8ACY6wNR9OcHTcD3zvZnixCqb91d/KpxckzEb4
jqgpLhpNphShJR5wnsfyk+cg6qA/Fx6TKX5GPiRhNyyFeUdfkpUDHBNQ60vBjXsDVfVZhCd7RMoH
3PYkgP2R6T0aYFitxufCmg+r2Hunf0Rcma6VO+Zz4N/PWSHdiIOzbUvqx4S2AOYq2LXr+YHd7ab3
cnHBQPDkGBrH3JV8iU/utZfImhn0US3VPaDu2aq9OKFjH9HeOe9omHLpzIlY5ERUvMqMW6prQDxQ
qL+oB+bG20Ykp4eyDoHM5iCqyeCBbkO6WWr4mwV/bgxsv/MgEcZ2C726dc7LDEO12Xyo90TAapA3
oq0Ok76NrIwuy6A8XJCOGzPeXkgpl2R5G5Pmyk/Ey5NPQMd+6XDBImPLo88Dj5h5Xkdw1c3Y1+2D
Ez513pGgRVel4Ce/ow8ZHQZFguHd1XDF1SdstL9uUD5kPSqrLClCWMSInWAexlL7iNjkczms5TDk
xMl8RpKThGASaVJ08YysB+jzFp9yLoF6evIYdkYrX4AbGe5n+24pxNahpCiPb1OyBhqeI4QgxJXS
zKDp28LAWbnjIGWWYGi49O4grZZQdHmDohF4u80q3sjiMfD6wox5BmoR53NGYsNWsjkERO6/hm7J
86l0JdjKrIb08dilqX+mpGEcwD/QiMInyiiqoQFM1Y7Eo/1ko1rFewQ9Jjj3AEkhzl0GZFiCWPh6
hlXg0vcHmK4R2SVotyZkjTYvzgn5v9WfdiSHN6N97LLAXO7D32K/1kVp9JTeda16bvZhAeWZrGtC
jXK094H3SH4yL4fieXpwKBvhy84ukXU4QoEKmjTA7nJkQs6g6RU79JhU3CT2M2eWB2QEihSQAOZI
DP+VLTQKkfTDjclhHM7LFM7+wWNRgAyRAA57rmtqyASrpAUdOsIvqfwaFdrCt9XSacYoO6a72Eu3
G2tFBirUlGjN7piBvyE3Xt45kS3SiaxcnxIiTGx41cSFMonpYL2k5yYtxno02+1JN3BpdP7CovwU
XV6h39gFsZDCLBS0ZmFlwfU1Hk86Ez3clcsimxyWgDHQ8mVyN1iq7nxUs8+3VkanIcPJS7ySyj5t
UoC+E+aWPQpO+jm5OEJ7M64G02E/OdmYtAUZcajsgugUfBVyO3UelMQIXuV3xR70MU4QRPm9UO5K
mZYIJGs28dNIRVhRcXXkyKijU9DNTkl3Hjw2/A7xzEYnN+3Qm+y3uxizORWmxnkZ5op8VHgsvAWW
OUK4shCKictaNz1qTlxnrpAER7R8KqDa7qWhOg3VqiwekIlgrW6oq049XJyT9LYLJaiCbToAUm30
7cMnqW3wzejzZQsLde6eTtmezcX3MgO4q8jd4ewP+xoST3WDfZ0OL03KTz3dpk6Mi6sjrznVAbTU
XfDgVoH6DHLxGjaQhAfzhGu6ZNLq1fm1rK/Ygmg4Rf5lTqxqnt4SwaBJac/9uCbZDOX4aKOoMS/6
hNrJDmKdp0591ZSVsOKJ8q6p7jM7DD+6h+99yTYTMCA4a7vi6eTklb5Yr+QMSOugS7/XSIaXT9eC
9pKS57/N8d9i77XhWGOlUatU+/j/FboprEm40f/jCTegdfH2T9+HsU3pU3ljzZMJEd3L3gKrG3/x
W5nZSSiNKL3JXdvW9wsBsTGXYj3EqDR+xQifuau4/ipjLxLzr5D9/Qc0CR0lSyuD+is7Du+RVEr0
Wwoh6fycgEyXxIL194qJMYLoTWZ2SndKZXcAEK0gGd+0qGG9yskHFX1ZxtA7UUOs1UpiZP4QKlNi
lJA/DtLn3QU3lVaTblSJHeJGruDGSPN2H+pbOwK4W76WKa/lRWwGA91DiGnPJlT6fUjAiR9RxmaT
v6McnDML6fV328oVIadCDdCVx5Gdck78ZBBJ6hA0bihaxgcSMxAW2gFQeRhjKTcR+3rsW8urWRRk
ofMJ+AtlnzQUBfZAXs0ngs77lNvw48KNCjNx6jdfZ7I4pGq7epVS3eYzcG+Z+Py5Un5rwmYnQyUq
3P+AoslkgrS/8h+KrjwxxIc0HJqQH3BMCYdRhqTS9Wiy0Urt7KtpFYc8mqrR5RyewbGCLplPvNjH
tlPHlHiTa+MTMdX7jdB1HIyPlF313t0ZRSSmta0GVtsN1cmW9DA4UjdqRBzad6ZbctVg3rInIqGQ
4xjtbuAwu6+ACP0h+6IQk6Ce2VBCQ2zpLSOJjMlR9g/NZ9KK9VzXBxZtYYEh6PZ96+HaQe/tU16x
06ANZtcG3U7iz/8hNu6/5BpwRkldJvv90OCMLlwvAW3b/RD1I5A1KnaWGsZdDkRokj505G9MyxHs
PkRTIVzFDwsmq2TDrlHHcIiD07+dPC1B951pdrGvea3vbUk8lpmwt0nILrFwOcZa9kv9Y35YOWzs
C5GxkI3TcPJ2+rDRUBVWKkiMyQLwlfVdPZPl0gg1jLaLTo/ewMsEjXfVM8Ni8utMn7bipdg/eLF4
JTT4TJpLxokmzrxXgZPmhm1MRxeW4/T0BK3ELB7bXTfQayl++TF1iEsxNCwHnOr81qZBE7uDRrxY
j9/5i/Fc1Q16dTmVgRmb774KlEVwmqhMUiv4M/7W0kpytpbr8eiqNEGGVdhsrrFS5qHV0c3yDv5H
e5QCYLY9//fXDqWJjGu4OFq3RtGuzTlQAoCrHDOrPg6yNajPvEg+yZ81m8+uuh+GOVFf1/X7v7C2
klcUX/lA4XxUnPV4ezSkKD+87ogv/1pNG/u7uRbGMoqmEpf7sF2UpYi5nBqziIuefbzjmqSzcJwo
N7NPwVvesvNbubBbzNucCECURDwfnzdQl6Kb2KCa2txMlyHifE9Fvlb2NN2FVrQ1m5a+jsiZGMSQ
xyegz/ei1uR2IQ+HK0azKfThVSa9KYj9yMq0t+u7TuxjWeuMiuMBpDFhvGtK1Kq1a5Sk49Vynpcx
Jz6zFIUQOOufMJLYMhQuWAOrauzovMx5WiGYjSXs8zV1iq52ht3dtRFlLlRyCkJM+FTfXFYbY65h
fTT9RahfIlaNQmForrpu2N4ysIMa4dT2Z6f/b/GnPyD4nIL192c85KUdY8LrnvzLmnRDpOC8riaR
sXX0SuSO7F/lW0IaJlpF2fjHLiQrhd0jsIQJnfHRTeTA78WlUdhfd81ztYRCqZZ0DepMcufbEOE7
PVJQl217NYAvfyRQSdh+cX6+xgI03CdNstk9QxjahM+58m5YOnP9p5diUII/BWX971weu58jRvZ+
33bfFRtfBzI46KK5MFNR0dnBBnwo6pe/2i4buQY5ugLfwrev0BN3ChsQ0yrTb8XbgVHfabuVu2tb
VuRxk6JddQxrjBt1aDBlDDQtk+JgzVgypT60XG7XvHcWHQKEuKnTJTsydHeWZpddjEsQ+DrBzIip
BRhNcvUXutQj+Psp+ZpTjJ2SI9WxFjI9YsU2+dIqryVSKpQcg5PPcXG6wIRmBDknEqmn/ytebKnN
JO5TrOCElWgz2i8j255x21ObVo+3Q8qrp1Jd+F72LX6edFo8vy/24Z9S2ySdO6yQjSdHkjLJwsFY
zRoi1a4+bbz0bd2tE6qM9yKkH+JESna2TqjJYDZWo13QuauLT1/1vnVmYGCQcpQ0D7l4m+/zecNa
I0v+ZqhYnRZLBFtnCoFp+RUm63/NYjyR6h8CjF2dgBHLHnwPTsriW41IpJhXpmjxZd9VT8yY8yHE
8OJExfrK0A+3+qtni8TpoaiAuhBJyoOZwp9Lkf2Cm4Jn+16+OmHUhjqAcJqYcICi8/OC7XOKz+li
GkCigzWwm3VnGjptKwEd0TE2zVOY+9DNKjTB5v12PED3m2yQZpbkRxdwDCW+cyMGh1FapN8KpOkz
12bfsjAMYeMfrsMq+LUlmk2oHH/GmuW0XZBjqOKAuRXHgyW6A1dImhepfaUpQJXGrkNh+0Tkzkxv
YGYb0h8fuhT5uQ+MTG/TKPHoNafUWfo7l+zTpZ1PpOzpfdja2f0+pNNBLk2xjxziC+AGZV9fm6LN
nYGvgL68u/lsJKaaZgEomYU4J0nanmgoDIKHn9O6TKAXpZ/3K2sqi51HJKEqufmPFxcMyoFgByNf
32cQVq4LYwbRrRPa6leRvlCoHquheBvyNOC/lYvTY6HWTfv0HkhAphI1tq5caXdqIiTohShMbzSU
YZHTCYIL6kURYZyC7fLlf07/kVhJUCsa2k4CeBVMYqXTH3OUeYEfJMUugy70mGh0jb19w9La0Wc4
X4P4x6enrwrO2IiIgQBjFgE7zYCf/OIX6c+hXhemWexTdyJvFn1QKWGISsJAI8gBK4VfUhn1KEgp
iQ+SMiO/baim+wNgTE6kJopCQa/4GImG0kil8nhE5AHMPLoDr/u6lgyCXxHDbrdnGPlvAS9fQP3O
Ep3egDaht2bnR5qcYvYARHkkPbR4guOmV4skYo4yQc9wROusCmEDsb4XE6ysVngsSuv4m1LUtaGZ
pBdAQGDKj4Qj8T2irDahxZDGpxlfiwkcZlJX6EQ1KqT9pNZD1UUzxKqXc09ectHKOg+awHtMjeNj
3ciHtYRR6/EhGJx1PPQoNCm4LC8JCRZe31lDpURYYL4zkVvvHbco7o31E/LV8+l9aX7cSDO2EoPm
UkT2T1/X/UsLFkSWnIxnViVo1roWLBVlHGvqHXevIAKI2HYuD+I2UhH1H4RJK78X1pssJoxoJwks
TZIXCQrqyRjJMpqTD87N9oSUcp590HqPPs+pcrPo21jDYhhNqsZMt1Fbrnq+7qwHoKBJVGufIeU4
gKMPqw2RxHMK4eLIgUPsi4cYaf8JXRQo6LU2zPGUPtfk6iMqvPD1FRnUPvLvVUeUtnVCEcpvjwgq
Pw2Udl+BVg3J8jyVmEtuVT8ODEomxbMWEkjDxwGj/I0aaBFMghR0UeYfXCrIFIMkUI95E4DcxRk4
+Liu7CefiWU2PUVko/vBUE4Ck96lTJ+MkNBabtqhS+VRy4j1akHk3oUw1Sy0HXOUg95UGi+Wawnk
j2l6p1ZWWGIrY4eEzoXPJEtTC5hbTYuYtHTgEx4XJSftjUm7u4gECAvIYUrF250P8hVEfHgwvR56
bE2sa3DR9laq+QQeLBwgxt71fBmHM2jhFubfjfCdsuzPA0lRA0IRCj6SitHGCkgu6DJrE71/EfZZ
9hg3te/ezYlTdfZPdVpSr1tc/3RBehxjXgKVQrHT5Wk3gwbu+xHux82vZpLn98gDvMv/WtjinTaF
u5f5quokp4IpcKPihid/dyz8wsDyEEZHICpeZP3LJ95muIQSnsR+vwfz1tXf1cN/1vYCemc8evpG
SEQCrbCvCqq2achX5gGrgsL8tixH4eO0HJaiG2lE1Aqdqs/KdabsMjClPQqkJMcXBe4eSLac5d5e
O2vXgbIlE+P4zlnkO7TMciCeuyRR/o7QpqLV/+G6KT5b/3KOo7ovsGljW3O+7yKC3AOyWcdzkhaJ
uZzYhpEM7SM1//591onz6vrNv+uT8VF8ywoG5i2Q5cotumbVauUApZ2vYZwmL6zOnD7HzbPbEd9X
rH7u2ocYIbBoOk4tpjQNQt7o0R0AbSL9/oGEUXv9XjHuEh2psEFbzD84rlj8h/9/uDikEz9MeWZC
Ohb1PfdkhyrEOkJDmyDvYk5NVsQzyGTU/zam4ecpVoyVd9xdey8CE2b8QdR+8G9grtE9NGs6XNAy
EYFJooDY6s3lV2wEGOPcmfzdsPosavvFC7BlEuZWL7fFDCbxSG0CpsXOJqKpn9lM0xy8nnWEztwz
SneqD3Aa67VDIr2dxggN7AgaM9xvFhWXvhpZ70UrXuZH/MGjfJ5aXexch+S89O6DYH33QVLc4caX
oUeowWYbqV1B90KATHDLSYmcBr9Q4LQ/Qob5wGqrEaRKW0GuCE1VuZ+nkwQr5RA1Q04Nxne7ZsCV
SHhhlF38ppqog956sHnhrq8zlQiDuJk6NslcoEZ4Ds4HT793SnfqMyo5Qq0fAxvxNe/gi15SH/I5
gazYozn4vhJCTuTrmDg8nRPtvrMf4R379wZR+Ht90wFMiFMIbOH5DpF5TkRzcmEqn3ZktA6R5JuL
JDRHKEWPEiBWC7zXbZ508atIjxJOfQbEVy1U/EmHLCBIeJwA4SjyPSuJlyd22vsmIHZtoLHNBOyA
xXUAepyytpdMhnT4lWaprxxBA/5B4lXvLvxb6AYhx3laxzUQ4ia9GScg9RJ2QyTMFOArhUQcYGtP
rm5VmSzec1zmky/hVbmBvKQQzvkj8fBVk8qK8CY6a8soCFQaG5lURcVvS/Vg7+9gXxvv1RFsTfiw
sj7PlWwbcUfE6eNoj599qfPBYJZy/lFLOboAXUjueKrTqw/vaotuvQ9Gnlqv9GyiYh7B9oMZpW4y
JRGtD65EEx/K9bhjxdcD+bdBranw4ptAXJlVfzlLPxpgFyRlrR6Whgeap0L5FjTx/9ZgypWLXx0U
5Cunun5jh3vzz+hUKy8L3FYPOH3tEXll0UWCE9Rlp0HDQ+Rd1Ypvq9JFABscdgzBdzDe3UOLcNul
lOwOII4hOv1Cms/ISaOfp5DGCbMleHUiGWgNFpN1vWzz76bwS92OIc+YIb0XF42f4EZkYofRWU0Z
FencuoDl1vFkhI05SM5nlRZuEHqsML58UXF+ENz8S+WCljM/8DSXHUBd9d26xa9iHO3pN13sgWtJ
ksAlgHCd/HiN6nOHVkxIlSiKZ+nSXa7v05wWQZCyhqGgQgeCzldcYALx9m61l/VY3JtyIIsLhjkR
Y27Hvtj9nQmHdDQGhn42KtG3EdNh22Aw9HHmfos5HJMmctrxYN2gwG0LRaeSnX3r49t9LXXkyHF9
V5+238XVjeEe8ShAxJnFHnhQXG9KHuuhOGZ9YP3JbTvMnxWAtNkLeq6nfjJ33PoPbTUjq+rg0k0Q
SYgWvSslPgSIAKa0k+JvIHL2MhNOdgh4HZB5vBOTRT/g6Tx28z4GKsO3e4PQ2wbCpBl9CCvdguhT
Xouo3a55J6KY8CQJbGfgf3vHTbApog19nTD7gaRN7I+DmpDLNJFGaPcVGnbPMlC1gcHlvOGm/a2d
DhDm7xhzOKIecA8qomzBktGCF4DCcqHT5YPQAgL1vmrgx2OYHURjKkRPzUbrARthdI/radCUnNoc
KfcRtSG7Oo/5KUGr/FnlqbgPquX9D+Ym1M3+RjPsrIBIN4PTI+3qphtAHzAIc7NVnFVhz0O6i4nm
bv4Y/UwwMhI3PoUcgTyXiCma3XeMUhNjxa+x7q1/NkNjk9PccUKl/FkMWdF2F24bh5YIP/hPfD8k
Dz6V5ZqB/+LeIelVX+53Y9OKU1lLcAYw6POtK0TfzTTBQPTKLO1L4M91tEmFJSW9rcjYLDfDSSVi
pTgx+vaKBVl0YozapV8h5zFjsOXAjuTqaQX5hBRmmCwTdsEdzmVR93jcYOjqNKIysOJlqRNf/C5D
UVDw2/05yMX7ou5SCTBxBWn46quKLykTGHhIpcpaIPTGHMiZIValh/jfdqxb34xnNQMVuRAqB+j+
JExbpt77v0X6bqgMW00gw0lTM3bEioFCiV9fR8sRcn+CHf9ZVPXIC7FKMUw0oEr4LpPgcc+G5JbA
FnuLOR0Q+OuJ5NLI2co7FBs9OrGBBbc+ZadYw5q2SZmpWnuWT6lFGHP9SCOaUq91PcK8nISGqScK
52/d+n/DPD3r/TYKAvfzA8GP4AFVEJnxb8ynNDTzVnoB+YAa5EKREYmeBDQdLDR3tFK2/zTJwsVS
AxJQs58zSMWYuN0Z60UB+j+tNGk4ByluqEejsKQhFU7iCvIMml2bkPNjEN/G7IISocRRndF9Cyiu
qo7ducx607dbF8WsDuKMf7lgQycRXVnQT2GweZtxuLeb4zATFT0k0rUgG5El4glJ/cQw1Zg7mB4C
He8KGam12KVjHNZbXtr8QhVuXTQsoWMpwg4/XSxguVWhPcRCy2GKZp0/s4VinJ0BcNKCVS2W4f6j
SuIvrhYAfAyQQ5cIaBYeP4ZaqLJCGz5ca9yuhHdrsvyozNY34w2dkBW14Nk29cYNmIdI6s7kigXN
VVKZcWF4mdQSKPie/tnJX/Awr3f0Pc+uImTEwZBVblVYh3a3ifZz1aVCeQxJ7R19pYxEsTJySC9k
mOxsgN4nWRFtDwkwPIhSpgmVRAae3LB5EAy/L7ldwVR++y3kO6ylWBMbzhryMomdbxtwApV9X9na
G9macnofhxGki9IzwYuLZ6vPvSaV+u50Fu7V08EEmUhpYrfSVo8UTsNQ4KOw2kiIlbT7iHfHAdc+
/fuQnm84SXQwJzRhWcKoTIwGj8rKkYHxzt1IOHiL0gupAR9sbqhweWAboS2Iyi4sOljKV2t9eKTa
ohFWUvVpwPs6GH6vxSIHJD8n0/BNvZuQaadE4Wffg+WR4751GUqixpPaxA+P7y6MuEOI9PF30KL+
Edl1d0rCn6cNmTYoWPCbVzOKQ9MIlAlUmeMYhJuUp7QzOyxBGnHyAIhiMfc3kZfItSUx4z1RoKi+
d3jo+vwA/AmNMgXiK9qB02MJmCrs99PxAElwwu8KVtHjtFCWOPaecAuMTRmvoCnKoO7KrnDLabdV
IggUVnlcquNsThqQHC/idZY8yGa0Xix17/mk/Axt3Xe+Ze2/a6tccmjDTPYxUH1s6N/T8jYyyU93
Brsc50ITptS1bGBTv0VgTy+T6lALyyoLTJn362j0/DGI9jwpbv14wT54wT8Ok7UEakuGsnb+z9CQ
jTWR3PrmlkyOivDY0/kh3nl8FWs1cOatIjRHyirhx9UeVWxv1cOe2a2io+09+c0E2WM8JhLHwcag
8/FNWX9l2N/MRk+5W27V06sao6uMxBktVplaeQ/7F32wy3X2aROFqchBh6amhm9wNuOssdNvy17z
MyQd8rcb+nP1dEAoW8aWjXsHKHl/nk3SbzUC9mDEeVhwCvJI5saHCXrb1CBp7VgITdr7qlz1MF0z
R7hQvJmS9t9Sbx45lHuurKaaOtiGtw2ZwnS9Ac8lfX4pHFaN+cTmI5wAO3jSg37sVQNgM4fgTM7B
yusxlEFD/pt6MM7ZVsvMveTXieU5VSDuS2JrTb55V/bCHy9dQE3UV1KALtuPQ+aNi1tARLjwG2vB
MKCn8HIMGn9AZF73nyCm8DejEarOc7cJr7UfOl5pyOY65fEoWZtGfTpD/MAwlooCypYUO30JAXsd
daG9D22LyNpLJbNXgF3jA2W5PEO1URrNQfosTLeJqMioTvl6ddCnzU2CZYw7I4phQtGwUovVkXf7
RVsNros5uH9O3QmIwEKiQMSo8lTNISRGxIvzczaEmkvO8EKeCCxR54UKggwCSPfLlKXsLXFGjALw
UH/SkPKA+H/iUm7VQrQCsCnXB918F6VYmtWW00d8YULNZXB/DCjW7nkkq3ipqtOXPAoqCnop27El
wza1hR40qv7gpGoykpvVAQcKVeO6HSa+sqLuOp4a0Q3hCj7FpQ72ygj3m+YHbFPGNQfKlsQ6SLct
8pS4h069sAQN6bAj6V9o2gAln6A1VPommLW2DsB5VLuNGv38w6jqPLKRwKT+NRo1lSTltWrLDlfi
HG+XnZk2UN0gPhQMNa1gZxMjTfb49GuokbrwYTQp6XBT8XY7Z4bdLrD/hLxblF3OvwR0RyZMb3Al
R/tSH4PrRD5im5iuhW08ENorXGHcqKchfMxuMRkKk8x5jsIzdezBHmhTwzRouJINYsiXKGP9qbo8
DnSPFgTqfrQXms+FGbH6arfy/dolimooMzIkzZSa4xeBSfPBuWnCiVL8kb/fadIsaJWLqIKAFmL7
dFIYsRF5HDQIAwyo3RpMfrQrp+JIsv5QB/bE8jsVVK1zZFs2oJVzQiaPoG+M0eiqHyjWOWYP6A8D
CaiHsSHAewQdea4bic+VfIsVtevhe4hn7Dg5MbTlBteSc7B3TdXH1xxHIbsi3o0podUQSVC/7PR7
uMOpSKIa1GWmI3R3gZi1Am6wkYEe5+b488Wfs5vIzOrRdVsfgvPVb2FlqUZ2B7VlHY58UuOoACPn
WM1kNrfPp+pgybwgaBOkRR/IC9g20cQA66Zd2qzcI12U1sAJ6odp4eB69kNfgqtVwPUsn7awUggC
P/qNOtvGNlO3vBSgRdtV4tWZAoA3pai2nOSjXq/B6G1ICJnryllKzlrcM3KAHFUNYs1QiDDPqAj8
HOKcysW6Q+V/dTHgp7xr1v3qf8n++khkAvPbTO7W2T6jO/oBaTUarChBFEjKiOdp/TZ30nFtT4AH
9MlDbNK4gFSmXnQCYga8x+7665OZ/2fzkGr7qFzwh42fjyfdBrRj4+3h2utmkX1RMTbc1etx0T0f
nWEBf0YJIZro5FpmcmmB22j2n/dDik5ExHv15qtfdxU47YR6GHIx2HQAQIVYxh0efZDlglDnHi0i
dw9NmT29pqyxJu6vOc+c8dKzf1c/ek/cEkTOt2v8AZVgBWzs7mgSfc2Ke/F2wldsFf+UkEcNYwsG
1NA8S/uVlXQRWzWiM4EO4gVjo05t1C5ArYHvUr/ENRfbGkR/QO+3d/7A4jhiNiOTlBW0Li93zuNX
ctzcPfIPTCwtTvOJKbPhg5gOt5ykq2dCbEnOYIJgN6L914eQBdKzdc03mnPtwoGeUu74C5IiCBFT
/0wQFEK3CK2msLeTjUJosjf9vtnCmISROKXWIdu+4yH/Jw9t26LC2V5hwVTRyyqt6JSqCHHyRtC+
OevAVR3cKEMX/Lotf+VD7BD8U6wnF7X/PWAY4zSYKwjS264EzLABt7we69F9zlw8BNclDmqyW2re
BZI4CMSdjluKjc08vBkKNCSxwDoREZBDe3+PiyYbyxFfNRHSV3Y5MrJ3iBG7Fed5KEfvCaCImXft
ThE/0E2S6yDhvx3v4lWqVp2n1Dqk0J+2Sk2CFMU3H7jKUPEmco76dvGkvP3LEjMFlQCFHWV+uTFO
pxpvLa+G8hAsst2sC04jUPptdrABO0wPEu7pbfhVTfHrg64Vk4M5NB15JXHFuAl7wHqkQizUlnZ4
BADYwo6F56SjdUoqj/La9Trnrj046qJrssnwHsDnHv5p85h3+bcvVcdgY3Ql/TNT4EgV9Tk4M5Hl
35Ody7DokITcKaczdaSktNPiZdrqvJzKjfPFlgGwHe1M1Um3+0i2j9x3KmznpRuMbr9tIi3bCbHl
htr30Bsi3mMEkyuyHPYWxSql/A2DgZItO5frgdjKPkt1cGwYoYsfVuE7Lwj72KMUjv5/Y+b7mdxD
EIFfpV0sDJ75wJeeYulbsQ6gDGIBcCVmcE2Y4ArIkEDuD4nv/xw0GAJT99dSA6xryZ/J2g/PZiXX
K+vZz+frdDUnTBcpKFyoP/8KPHacuR0Ub40kOxgj95R5HeCU61MJKsteO93V52Ckgf5/svVuFo9u
fjsUbkX3hDUYZrrygBniiGNE0jCklebaqsx7Zet8rHTq6pTzA2wTcTfZhTITEOFthGgaG6FWRWZ2
I2O8FrfGkd7wQ86PxvpI3HEq2K8I5dJTIw+9AJ/EHeNrSy9dtwl8zu4N/nL3vpUd+3yGpvWJ//s1
Kz9LZTtPRe/6If06MtypcRCdp3N5UORQNzUVZKeiSHVvAgzWv4D/28qZzVj9ADMlHoGC8aWo3Wli
uqiCFpX1+0QpaNgJ02HaFxp6B+S1uBlLXDyzk/zo+vnbE1uYGL7PfFRzTJoYDWWJXC+twoz0UZ8d
2NTFzPyuO0mb6lDK2UjYNiMY2scWIad6KsS03I4gYJro+08ODwZs0Yzk+wGPLKZqrswvQV/NCtjB
zLUszR9jNVX4qIK+Qvv0wO83T/OFhYXKtHB0pWi+G4QstidzSGcSGs3pvRVsGQZefPxOn5xDC4U7
8LuEOl/KwWLBGExpPNnMdNWWAfkUMcCtqtDoRciDTWqYT2v6IIZvx+wQ8h+k5zfOMEYdyfmZVIM9
83Nf0Sqma7tSc8EUNkGkcguul6ky1XoG0VOf2r3tL53pC85iqX7Xc4+SN/XIN/vq1hJvqi6C1ieR
VTy1+S0O2WeDdO4EjgREVhehOakUkegpGzCazjPrziUSTkkRTmN+BOrwLcciRSIBNy90UazPsidm
wKZVXgRBrl2HFwJ1qZd0nBAVrL9MeBDb2/6HFf6cCnV+vpi7PWWBSDy/aLOd+8fzcYJ87IEOhmTY
pp/vM9aHLgllaKkEelxrvqit3aSJT9qXh6wZbqOP4QjfOS+TE/cLJVWQSIpBWQyIlCh0Duxa2EAo
cIJlAKSCtIVX+rOPX2FABBnXQu8JOQP1ckKAgYgtwr8siqzinbVA+0RQnLkF5Q6bBdSl7LORGstV
DII6MJjJEHzLmtQTubCuxRRmHoDVs7bH/PamH3100lE+C7cnpjh5TX7NUUc4p96aM5ptVgn2nRlF
IpcMOnDpnmGVOAqbaQcmUyzYt/CgfLyHS/t2esQGye2c52wN9ELcBkJyKbXMMI69T9D6zvKsuNBU
6hOLrTVN5A2OWgudxOAr1Rwp0b4YWwZ+haP2UB2Ip6Wp69NL5gbHmVwBgx3JZ6RlpBGRevQN+N++
idsOJtPwhQytG4s7FMh5CHSs1q1LZ7DCF1sJD9bai6uSu8o4a01AFl7HUdDzFAXndjCe3a5E734C
PE9x2HtImLZZiY1kQQx2QHqiwqGwA90Pn6Y+rsqLacGysJj8/5wqXhVjOpBTFwFt3n4DWIGtlI+p
jVhmigcuZkDyn7cy43WpnxyqBZNABcdsbwHH0IljIUSpOdk/UdqR1Gj+qnYFlMOo5hNOmUutXYXN
uLZHjHrm8cdvzJP455oBCLXBoaA65XgfaIIuhvEBPEy9/TlZtHk//QzHkLo1rTzE9oY9r6PFgKjo
Uv3oi7C4EtC91wfq6AkNdrDVY9/JAt2RBbete7pMCuyrRkGqzsqxT+PvVdM8HdnNHCWbMi75whFs
8jSAp+Hj27iq5QmFhUj7qFCgkC596jg/o2pAEoL5DEiJI9XUAn9y92A85e8WTOQqFVP7nnhhV7P0
omO7djvK2Fghrbue7mb9YHpoC/3crBThN4je1nrH7hYCf2Kq6Xmypt+MG+/yZW3ykGYW0BcRUJOC
6gq5xdPL/JsD2k62x0i/Lb9qZnBtSzGJvXeIBTfWs8dRd2dUTmTSAMlYHzieN5Wua3/RmWVig+bb
/KOKVBwwDS+sfrjjB84KAPt4LRp4E++ild1Ot/jycdC/MvikoPXwdkqHAF1S4jG8CsTL4oW4fMOu
agT6TZo3T1xxiY0ZqxcsL5bU0A5GDyeawnoBakQncZAV1C2Wfs9tkzMXkFM3qtNEP1yy2bZ93sdK
IabH+nlAmsHoJd57YGq3v51+IdZzHhX5tbX8n4cNIk3uz285sJZeoDCoqAchZMEYem9XzEQmJfkI
H7/0LL2d8CD8SDTcpo4g4EP1bP8jxGLTa06PACltu3Ek2CYETwqNyhaf4ioDa9ffIM5JF7U7eZG4
BDzEtV6WORLbVZu/iAsimlyt0NyrW3D3Vb9N1LJxLe7S7lqq011nfMwT1AR8muNWF5PkmEs2a77u
WsE886BnZyU7DrDS0v+C8yZhQGOA7QKdHLqdDp+eRaELMCxQAfoeo8KCgqPfH4X5ayfodm03NBwD
L8GsMuMLHwMW93k7ihqvK5pJ0nAQu5p3fSx7LcDTx5QXKrf+yuhwnS4JcaxXDMBvnilxRjy+sJdD
LMsDtpRTQyHR1NXtMxAWcGuwcKjJLiq51k9YVcYUe7tSGsS51xmMaIgpJb+yddfVRj7Wv5w53Yk5
hDbxRnCSWSom/QX7x8U0SLp1bE6JpT3bd3vpKp3sdb9i+qp23puQGILv6pctzc8+A7Pwf6d9uWj7
fFKxlu7bRLyOoWuLttw/0FdRoL01/qgdRMIfbqtO1cXTGlB0BWHv7WGDzP0M8SIjS9a8KLgKCZR4
9rq+Bk8vkFIbpk90WQESsTw6jzscpsWkcz1J+/jqDnhiU6wcTdKuGYZdUPcJ6DbdF1nhk+K2aKYN
IjJs9cj2jCrr22ndL9XPXvpY2jkz+9c9uwDdyv8hBSyVTwWeuXlHQ1p5/ZRDWmeQWXQRP/f367/4
OR29Lo9AYBi3f2Hu1w3PhjeYa/Cy85L5uX2TlzSRMy49s2vcZ3ObgSu1ehMgOikRJGVeOuPCZr1Y
z6Tsyqnon2276AD3HZboDE6BzyiycZLSAJGcxKM3ZgWq0rd5sLs28/jvmfYeqOfioK7PREt0BiTm
khm1rsBPWiKO1Ho1JeSdBaNTNtmjlGZPa3ZQjnRSEwWnwAeIq7uUSUjmc+RySRDjojyla17T8JUM
hygmX44b8hknN3Ms7Rr0RrE8RI1lWAdHP7MDq4RN/Ug5yda0ODhUjAHXsIG89pvpFeKSpmJ2tj26
gZuy7+WAlnq7/HJk9e+MCVDKYvpI9EFi9pEiqgwJ1Mi6vvaGy99KlxpGERSNWe/5NMzOZdS7E8Pg
TbK6EqX737uQkL6RbjSMyb1/ejh6dNUQcHwiMAixrrdokqSei11eBzlP4Es2WGer+gMC3frdladR
fBZJak9g69BoSdtudlGyFk1Z/wgRao7+87EM7+yoqHDlbB5A7RSHgqWRd6i9/3sW1Gl2e0KTXDdk
IqS9AWyrSQRWuSpUY30jjKboMUeNsPOQzg7aTmzIqwIGQ7wil34WPuEcecUhw1onsSyNsBAL4Ysp
YeQlUafF1ySKWsCnQ9VUsxrXjgHrEnHqKkbrszNlgxWs/HYqgKG7X1qOTCL52EXwOBQM7ffa90aE
BcTyKKt082dmyjvb8vuOfn+OXWznFUaRpDtrOivBRrOWhy/HL8Jtb7NryjY/R63RIH4zoCT3uDEj
HKv//yI723Jym+BQpSuDNVhaOepfTLYsOhvLrXW5N5LxnBXzE4O4FKAkhXRZ8T19WbKfqLHAXGjR
Lz7KssdPAjDYm89en6pB4R8Bs2g5d1GHQc6sPCFV0vptYXIU1PXBdosfzsLncZf3tmWx5jGIEybI
EMkVMu/wpO63QkFfuxHg2Ng/LuY+ah63ixotM40CCKv7AsrNzmzHP7yTQuZ2pYlVOc7C68EyxNEG
+yo2FmhuNV01TXuW++TC+fmG+t5d0g+ycb2uRCvH88und0NJEBWn4s5hLCom0nuZ48YYMM9lmrKA
rQJiJ0c24KVaT09P56PL/SBiqjtDyTmTuex2fZZUrHFGRehTxlPR6gN6V6OJM/JaQBHPJqANIBSc
qI/yzsopjzAk+akpew3drgt+fxKzGauQPZCEzCAXmWvIpou8ebe5673osTzUlOSpyQL2mul8tDvU
CpVHfcF6h1ohAn0Q1K9XNXR531wDz2ZDeX1evCeygFsK4Iah2sNzle0fgK7UFkrTmOLs5rrA4VpS
DTs/0vDk/+gOOXSsuvKXUT+2laV5cq31A+y3Hqv8cA0BZeCINuGB8K025GidRr4nYrtY02i5LsEO
gNl/E0OvT9MFtKNqSCfe1+thpl7ZWovnJ1UTiEUY30oYp2Z5dN5SYVc9Nb9HdCE8ZAG8aLcmWbt4
Lm3HOVs803pKeNOBWk3fpl8Bm33EKsy12fGTek9rB2VnWND+Aq6X4eDzX4MHLszoqNLuwdjokZRz
uv6T+UeTuDrc9BKeZmsQlg2K/Aehjlli3Otpvo1h9asBPc9p0jNotIBT2ik5MFAnKjiqBQCubHeJ
Nk6ssUywGZIz5ihtKw1lnDEJZezSqf7QzcQ5K3ogW+B6lQKtKMHkQMa7SXQvSJq7RFG7r3arKXmR
Gh6QP/7Kl2eLH/RtB8uO7uUGPKBjzWMDDHfWrOaUz8490HzSoS+2AJs7C12coxLBRKdjStiHO9js
0AQZ+WV9Zvpb2TZ/FD+vYtje2fonC65QMWhfSCSKDfKS8YKYeOFrasjSSUDGWs1gm0oL4waNobOL
ki0T7etjJ7Gx0of8/VmBxDzO8r8+wAw3ow8BrQNnzaNldxgSzl9NwmRYYPmeGY2QedQXjXz5NfQz
5FJERRE5Ero5hTkHi5A0F775L/T2/fso0pnTegVa0hE3yXEbiHiksobBu7NNj4dgXj8ony+LLFbz
uAmea/MUB7U2s7hsZWH5jDKBIi0cuqBTVM+uX2gEHvNWQUkVs7x8RtnEh368eZoyHLx4YcTdYvUU
nZDBUE1WVZYdiCxtP2DVoXs4R1L4F45vmTiZA0E6SMJUlCddqLNGxWBTipHX11m9Mc/P6jLNFuWa
j4EMwYQm1150anbjy9mLPPHZDrSLUZriSohqgA6ExLUms0DZD4DU1gDWYk7jRRc0pk7Bv+CrWh2n
LnNTPq3Sx7UFjFFS3VXI659V2bBomRI8jHCvTOwsUNbykUh+qROm/KtpkDf+n6HdTlr7FRZ6Lksx
HMbZuAxevz/lOZpJheyP83GF+p4RRsaIuHUEr1ZGf3+FLhuRTyY6ZswaQI624oQEt3afpSdTubX0
CMLHCMxbT53ubasNxxItYDttqYmC7DzWR+xkvRq/4lR7IvzV/WpZImIx6+h5pWEaeaEJ16EQzrgp
+vWGnXtolfnUNBMYTEsgsqstFwOPYRPWroD4N5YL6Y56vtX1nVcQk7GpYxrJClpo0Vkb9cMWG7+B
/ma+aUzLn+CNPNpu3x1ksqm9ORzTGoQe8qyYALYOOx800OIeGuOQUrZ3tVRgw29MOPdYnnLMO6km
EGmEoUjsz7MtcEk252lc+3ClwBETfwegxIW1rFoaSkvzqqGt5H1coeq6VnJutfGREEPEBXuxp1JF
fJRQGfQIc2Wpx1/sbrztx8IWbmWHV6ZTquKHS1I17zXbN4N9WSc2aDuK18jRP2wvbH8btG9AL4vH
yKC4nl2rUZnuiYU+1YWZmNYQ4jffCexqpX7ZCakDdkWnjArYx/HVtda2MWMno0ruf4ai4zJvJnTT
6VBJK1Z97YiNgwtrT6Ka3ucCMvLTE4YbFj+/tB3eJw1Gcv8afNZ3ZRBOQVJwsggMJTfYe2IwvzYo
8r4iTWwNzqAc/8d43qPQ7IjK5ppmkFFmdp75EVNchlrnQkLG1quBgiGfrcwCnbjExlz7mA6SedL2
JPDP+lVQfTwu6iehDJcvAWhmimJeFTrMH6E74HyCCWoiNA2Ke56kc/2UQ4uD0qc5bgnTkCo8Ey75
2t80XwQfjtk8sIGj92RY16HOWr/qMnOkDzHf7vVNdqUev1ZSaCCPpRa+Vz/gwRE4m61kCABCxs4u
ldwoc4NHToaByGJ7MwFFw4vI7eWaUAAHn5nIh5OxMhnoZYt+CSszDEdkECn1/nAiXkBzQVXlWg6n
82upoBt/5fC8dziW4+qc41zMWHdphSNTDWfdVwVP0zjuholMd/R2W22S0Z4pLsTFA6U7C1XNPeC9
n3fhUzyTZvQuuipoUVhyEUgtgn+kXkLwBVS0ANQ9IwimmVP5zzo44EyQtpjNJgvEw90Tjl8kzySN
ajqNZApHpMHTCSsR0vxON1PSEF5+X49XJ4RAykUYfSfjd5ahcTM8covZnzFKAsN9QRFKHarnSbzY
/qvGAWTD3kvinnamGCXGw5anCs7U60kFJ5lXTSsfR0WvpDY0QztnCc9Vsgm+0wfnCHnLFkzgfgZG
G2juhHirlGFsJJWkpC3fF+N7M/56IcSftuc3S3yRH+1sgUUKBQRvalF/W03AhbP4xlg1Dm6T0Suu
Ws7Ptg7kuX4o5t2JaFryyqPWmKktA0DL+0/hfYQ4NCFl8LBGjB82B7/Ih2V6rRtFcwXBnjiDYbCq
ub2gqkDoSEM/rcO66HJ9ocJHOPqFQPxQ7AnakNXuvxgRRg9yzpi++06aQelGiACtpAK/lKEu1lU7
et/5fHBBsVuLEC7hJYqnS4Il855Cay2DYpeWYbdut5Zz27/r2PadqC2MdoNy3aNR3HAdJwY8sJG6
sJs07RYNP2MNg5Nvaiv/KGwnC9fMMu1via4F8TPDTnC99sE27GnKiPudnNChwv2LBa/XLv2PLeQ+
q/pBubUXYaLEWpHe6Cm9fUM3g833jgOjqGLd20Rm9t6OROOFuR0ZbcHvbi2rjK+ZIU8wgNaBfNbF
1D5630Wn+wn0HBn0FeqzDfNEkWkSmNwoVsQYtV2bKZCHCFkvKb5U7kRJz6+lzgMF6FWMVcuRvvBC
bQGDzbx9MstAGgFWDGs05Id4oVt/GzCrW+zNCKMb07YckPfjleLz1SjMcHufuWke+efzKDRxPHtL
pRU4CKsWbNgml9Enp0MwHld53IGHg/ecyQuXph0M7uCEqUX1v+JMX2yqQhSOANr4oHiWwP+wJpAb
Ja1dZRrFmFm2akoLtDjMnGOFZRdmYYh5Xk+fnXfYau8T69W+NmLSXNK4GZ4R6XemAi1lI5whvqZ/
LgRho2zWmZA4a4VQVIBWtkAsumpBntSj5oV5dfp0HhADj8e5/gHJ5N0k6IPtTjmpygiH7D5VWU/l
TynYxrra8dOyZ/sWJe5BiuhRYIl26hYajvykgvjkQlE1tXsfGrtkoLCZUqKwYp+ShpJNPxFQWv3I
+VwV2F859LFeC+l3pHPGHGmkZvs1Vd7L//dwysC2CcPUfYdz1BM9SgrsLZFWAjnWqwRnoJKBvNp2
xgkkcnBWrfOjFmIi/Wxx0yscDNJPbGPLWu1rH6zBQqiackUDOJRokH1ZkwAlERJ3EtDL3yBXUbsT
R3ubGZH38lR4KOe69wdXcF4zqktYBh5aFYXtoLXtDdum1hzHZ7xwZgzRvgEC/DQqhMSKEWgKV/65
Vent3Qg52QFOrdBbuVHBbmoSZhqmalAJNg+JViM0cEK5rYyTjQBL+/GwsCkadRCh8M1ReOPHyAWt
S3e7IUfCy0Ot/C9zAYK6Eht/57MktCb7DGmdf5B05Cv9Pac0pVaoxEqHIdOFY3HHWfTAcVjMg2LG
ijRNnlC6000FzybJ/y77dEjhygb/BNPWaEzUZGCIvOEXRwa2Yx1uP/bQrnsE6S+pSIj7KXtmfd50
GdYVZaCojf9rxBSmZYLc7R4QhxX5yjrYzuyzDAghLkZ8h7stl1WWs2kNljr4C0Rnl/ELulNqA8qJ
/u14mfzKKVd8kzZ09ts+sMFW/ZPFzdTWEGyuBHkxhmh8aKKr3d+OU8jLTdJ9473vj4NmTtsXR8uL
l9SgQvZvfLfj/NOfHUEYv17FwUBBHNsN0ICSZy1tMmxBK9n5CtpIXTqP73D1orcjEIHmMF8ZUeSQ
ctdhO1WmP6YTw73UuC9zFeIOT4bmvprJ+eqxSAciLLFqpUTKKtMbdGnHNe53lgD5nbQRml12mDs3
7B1TEr3fM8EOlQhK9tKZA1uBPzN/WUjo/HQwsK9Rg0YuSJU6dGw7JVsXng+UV39eV+j9l4KjkFYC
XqY52bRe301PCVwLsSn8lyI8q4De7hGm0x+DVMAQpq0GuYYYBKmi/qL7t/KfsfyU+uTj3zp6QkcB
hlBigqxblZtRbWLI9ryCop5HddJUq6hG3ZT4ReuvT+XGa7UGuOkiJDXGFelNdNR2rnxiUNjm1VS8
r7SDDh30Li2B0cwe66VLzaQGrS1LY27lSGzchRyg7EusqVEkTP9bTk1RHVcy11d3Zi6BcBrS68ZX
HhZd6T5rsc2ovpsgv76DFrwVJ9xRUKgz/3iSa35c8PNfImwNJWzhBvDmUr+2kSZ6zGLMYkVHRF0n
r8dRdQNJL6RMmn13vEuGAA3SAu2X33iT6hbRtlDO62SlVhSBHNUgYSd5bslRkq0YvUzZiKYbzX3D
eE/u8LUVI3sxrT5woa2M4HmwNwkYjRkxPcsDIuRybhaesWpxciBtICvzdKLAltjWcWCSnNSbJhjk
JUYELOuP9117fbyRE8p0cCIiAvRXEUC0QQ0XQ59tOs6sk/AhxKOLmqEdbSG1unIK0q41820S79xz
cslB3H4ZfatiAlVxbDX6uBJQ7NW4GXfSTnErf1CcQqjVqt4q3+ewCEtyUHP6whPOF5rgaC5kjsWI
qYzIIv1LhD38ZfwWb7lr/hON4VFKeaFAGpMqOTFrsJ00fcoF40C34opwyBnMV9ERBL/4dXfajekB
atOGp3mvZnCv4Rac6vPmdN/o38muzuobUmbdZTxMVQMeg4JWgxru1MLKNHgU78m9zeyG7GNPPQZH
FwT2RmdZfq0YzlecY5XN38eUMMPzw9P/gILHzgWVz1ULqYAoS30YifokDCJ61QMFl8GmcJyKtUEY
cYKTvnj2xZYFJhKdBcDkQolYuWK160kgxboqpM9JV7dmSLBp8f1tU+4wBIBfcNZOx54HrRUYvbpE
mvHL36zEpCuNdnu70jqpTvdmnoAZsk6UPMioZ3JcJvJx60OH7xRPwwfcCZGUxx0rdpaPVQDNAmX1
Lf3+S6VwqAH8gWsMy3qogzzrd70KefTO0aqEfID9M12JFUPZsdD+C2wQZMCAWFiScFxcxI8YVsGw
d42udUMTcBQjhqxvcJGybykZy9pP7QRd/cQmZchdM8s5/OEq7+srarTp+6OpgeRG+jYLnpM2cW+c
Ff2dVNtLkA6Fys63MJngGnTv95pOdcqRSoU77pbXhYVI5p+oLCgVGpL3EpiBBPxOKM7YfdSKdLdX
fnH93BaaJrhvj/n1Zkd6rIiC5XVm35Kll3VfVbrcxFRkoYdyNzg2X68q7BTyILQKoA6XncpMvX0t
f+dgkpxQvCAfisb+Mj2IRueOQZR4hKhEh9gxZGq3YzUOV/IKLLmrgESWddz5ZSjUxqBZcixl3nro
Fe6z+gn6yT6b8BAh0opUrOXbEfTb/IP7cljrj97XBf3T9HBfp3shcCbTFkUs1tI4r5n5A2Fs12YB
PDLCRNCjGMwDlBDqEx3cMbb0wv4+ALlcr3GfEu+fDinEn7Bg89lTOEF7ZyySZX9p25kDWWD+voMO
Cpa/44qqJkuHa2WMoLCwxtEJnI54TpBZv+3L58WeBiLKlUNtf5wIjjfCD6ZEGHTVd85EqDrhdjNO
jnBvyy5w+UfoUcv9BqlKY+9nyl6DLe3a8CkJSY24X38/q0UZrij9Yzt3LsmURjgXP360PiiZ4ucD
IPjN95qW2SkGfTbuuykjBeQkTnpjthJArSwmkQxqEOob178/WFYjOR8pzqHascqCbQR5cHMB/Sim
fpIGb5mHaA+TSm+04W/qCIfUV2qV3ZYuyRHzkNkunY5OHnL/T6uxe5WNi20GzSowsNaiYffv7jOs
IxhgbldGWqaIAqIGufVHE83eSUu5PC5iqvojJXXBGjkWuS8piq5DiXybxSuvYk3/eRa1gB4Rq4Wg
NjDGR1KtDST978lQRXxXWW3Ko57jfZXfXgCVJVP+9rtLyWX+NiIvjVcgUc3do+kc9lsGVXabTQb6
9YVbvVXlHgDAVRF8A9H5hoV8ak1eKFxfl7q9MTDVbhOEIL1z+dk926ok/FGoLyGqTuzJ4wPyhuzC
cMPAZRNS2v0bxk/lADJCtr4cd4PNXroa73GEBqEtTC9KxA0Vk+IQiRmIZ0QnlUwuzKY/zp6y9qig
n92IRpHfDvmaQWR033dhu7oETDMvVSso1ysmlQa4Z78trTEE0bWYlwq1DCKhYZbPHrQOsDfzYzOx
X8A3aU5vfo5QBH43dzHpu6T1LZ7AgHyVeNqyxivB6MyhE3poIHoaMfNt3Lc9mXcvL+6i5tLd7zgu
zqBJQTupMX6ve23sa914ysX4XechFARMaZtguAg+neah6p1IQ2CvZet7pJshS3wU9LRtHhvmRZlf
Amerhm+d6vTVtzDOGTB5g2ndMM60cGJ9d1+DX1emEpic66hpybjipnqIRk/ApujgeM6hdrrxVFU2
85mqdt6tEBjuoakxZHSDFZyXCPWJ0HVWLSY8ONcCExoUScNB37vF1ITOFUxD1zIEBv8Vt3KA6vb0
rxeCpIxlBs548B5VIemqcLUuAKRryd8UZCAG0eSAssW/PMPGCORH5aH0Jyx/8RZBkc9uMXw8CPD3
G9bgQTYWnEd8O1mhgz9v+tcfjKVPLHjr3ME5+MWSUM8oxcZiZWPQRThFv4f2Z83Uz3b9N+rR/Vbu
yXBQkehRx7KLtI8ID5MOOhNwvlNyOcdBGX4cQ294nqI2oUYN2LfYRxc0gfVdRpR/1T3KSNgj9CTT
xdt6bZOEAGCXA8SsG+wmU61nNmbq1BQZ68qzBr0rkmDYDRO5mIyn4nrmv0ucIKGRD+Ar0QhfhWBM
UwlLHLojVdw+UA/yzDWOBb2jzDC5/MkCcJhpg79nfiuZ/NLakk8vjYdOIbbhRU55n42/Z97erVgR
ysruA0MBERSdndj2kkIeNyvjctAznFm4GhynF837QOSaihNUWCnrXbRfZpfIT/QVTkc5Vv3FclL9
llwmqQRWdVXJdIz35HTVo1aEXlLDTsDNDvwCeLuoIMk4r4jurrEPRK1BQqzkK+RnA2yZn0r8dfVZ
u8MhbEhB77+KT2EIODAtGAY3epFLnM/G96LAnk+OB4dtMSm36SjmmBUi1q/nmNGMzyzz5FAobcB3
Ra4kiej8wpol9lMroUPDG1D+MXCxwjGPYiUjZaJfzcR5rXQskPqYC9HSoE4DkSr9ruUc05rmX3r9
qYKCkRIM35IdD8SB0/pQ1BaGUIJ9WBnu6Cckl+V5AauSNGUKfCwQ/LTPiFE7lGlK/t+UvpTSAmnT
EqGVYUM54uCusNEBWgZNt+lZimKeFZgBE08iAoGW5AWtlE9qvv6X8Ixit9ht6NSKwbjadk1KO8BY
UZVxeCOf1msU6UH/q5U9HFSUCwJU9g+nqf/gHdJK//cePhBqdNUjpvyEzqyAjQ+ZUJAumgFW8zhz
mau9u8U0NNgWgTLrcqglGUr9QWMMGDTbFyVA0kGC9zsH7xUeivZ+/QTnCGHAcyFcY4Pn8MZMhxUR
OYAxAMuMNoGxJwlhDkdDFGG9T6dz9b7caZ4+R1TMxQQcnhQiYLnuk/jmcRffoO+YuWb5uaNd3SNS
LsAdgQpCy9qvuWQfKSbBU27QMKgf9tAsWfPi2jPhemIaMYUTC4G37oPyrTknrtxuLHCxEswl6plQ
UpDETnwP6w01ZLbL1ulsyO1qNTT2m0Z754JA5tksGbj4VZC3aXkE8wfcZ7m5pEXWPxkd9oI3gG2z
kQzsTY8+lI1/1VwJjXv9j/n43kTAFEAUAXmAYPyAdH57xpvaALwkzKXVQWUC75Mp+GvM+pPw8LUH
DIzXzoW3Ohp8+DGotYcNzxT44X/vJJqwCjE+/PMHwWtIVmvJkEfEFGDPpUqL599fXBoakkh7oht3
vO4ELSSpUxU1KjUsE4XYijdqNjxfVAvvGN8oysoLVceZcifjSK5+Nw2WD0Fqn4A9O1ed4eGwR6HZ
K1j9FCm3VGitaReE1ILDM3Y9cndH+MUX2IoIOUu7tYdV2mOROtoylVtCOTW0LOiX2lxnK/Cqjwhz
g5BfEffq/WnALgs+ymxWrF0N+Qof0tGExOTX4N5fz6wo/WaZcJmNZGEQiHNnt0ghSXquxjqV8pFi
1/STefSlAJJZwVMRRSgYUDVMfdX2HFX+SUZhbb/w448/8IGLf/LamxHQV5qQ2JE6phVoHccIvQGO
RExa7lKEx+24kg729FnhNCiwBCQ3jqWBQH3LGWqMtsqBV+dFtI1qMxyGTFE6U6vYBNWRyCYtpZJw
yEX3k/a4c2VnzKE/YwL+UQe0F6n+LsyaY3z3lshDM60eMzUcur5kQlmZnqwuuZtTdPw8NxZ3BGJv
Wn7afAC6L1M72YPoKRbcvKFfy50rfm17GpYVnUx8vIf0ZLgGUpA5+3ZlcXLOusw2jp+S2KLn/Wfg
ILPLhZleocEziSCytbcIJksmsSG3ebKcJYcuSwD1uHpN2k61/ZLjL8N4W28vpfOMaV5bkYZxbDTg
WhuoPTsLOEgkEtYKXHI9ymVgw9X/AeP55yKgo9bXg0jlYw3fS/VIRHRq2eTgijcZEz4bOvG6AL+f
VRoPi9k4irX4PNo7p493QCqNajz2LNPnm2sa8Ex9axm+adt3aKXsQbYPfNG8TekNKDJvtYNokQZt
Qs+w25L4p9R55lrGbrDHtN2pJKxgraS5Jl74X1zEOZXRIvG3rm6oUhAn61sc0pyM4dogy2bWGdqI
8/KaXMAKiMJA5wMGBSkaz2MF92Ky5Ke0WOdvjfnrq2pTMeZSnpQeVdK8a9RdWWK8JgPWhUAY6/3Y
LFVvVlsEJeXiHRNBDurCfM0OsT88h1D8w8c0U9hNrCzPzPtdIljKqHiIlzd8rSZkkZHVEBuj8Qz/
ETY2HmU81U+BUFL84HHnHiO52blJcX0iTUKnJgEet3E3zWUUAzCDZlLIY7POVMeTfWhBUJ1idtBh
vGySGSKEMQ8YQ77wV/n0Q50sz2sDeykH0MRiOxZYSxmu6zoKeH0Q7gfuxHOfnCybCSn791xUS8q3
haAzDsydgYAYVs8qaMa9/mO6awkWFH2erH94z+c9PCa/fmpgnuH9tWl6Ladr01bV1PUCHICinQYS
pKuXHYvQnuicXbMr2cZAX5COi5vXYa5utKKs0aMuaqxrvDsKNChWDRx78Q3+FejFSS8D2vniABq9
BlOyrXV6uRAwJGYgxSsHquAdCvWqzhaYhlf4CRJczKuPAiG1todurwH9I72qOQZxo8Y31Uln2rOA
puwIOuqZxh8Qk4BvIgAnKOvvUthaxfLzr/sJ8/OM1FAPkhkQev+BEh/66bnamQknu0Ymw/osUiTX
LLUBnO+0IaOQ+/fQbs7MEdnHja0V/tuZS8gQH1CIbARFjHajADMAbkMJC07tmAZhAd2JBlcIj69k
gRn30HAas1j8hhQXnv7PNGtDfxTeuwSkHrrGOSj5HlfxwoYBps0Q7NjcPobQ1WE1PddKKhdrKlfk
8/RshlSVQhRRv7AoBXX1l6lUmdOF3ccozJDj+ADBZCLJV7lX7OgnVmm9rSEtm2/aHrtZQVYtkBTC
XgCC8rcfSjYuQjm+pGQYv0j+QrOsfTrw1JUDP+hEiYJlTmhEBucTerAtAeGtMQKKI2VlUtIVqEW+
w8YipodZh8JZB5fRHeUiLQdn6541J6h58GI8ivzp9kulIod6YFPSCMEFSsrqKdJFIDrdMkEyL+Qv
4sm9pjmIfKYPGY0HNgShkRR+xQ5HE9tuB1aippnycgKlue9Ab19ltMMe1dpVrk4doJhKyWuW7dFB
Lm+0jWHdFiINw9vIN9llozygMs2In62F0V4aOPv7p7YbLi99lXtuM+e98Ug371HX5OQbPt4cJy5F
NPo4QHr7CN8stoMssmi/O3fHdpMRzXTWdCO52FjPhl/dUQEbsmMe5U8l2EglTPuizX3kQHlbnpKu
XiB5A4EBdS2zy6ZcWuDoJYD01qmbZZWG6j1I2/xLE98qH4iGJgaLTueKwRj638MYFzlOxFCNY35L
FjEMUSYVyFgwdil39dWSnqLNdQGzlt/0DnXcZnk5YVZARa8SlNRFZDA1Vr8dIdPnHvM/2ZA8xYEH
JVeuo0Kh/OkbdMwvfFAeQZ8LlwK1jlZhYy3pnQT3iEbTlERPItk+rsz1jeEqPoNUIuqfgKwD9GHu
FZHoigCOxSSQp2rYbuu8oS72MLAr5rjDAZ5HzyKpxvx+R2rOB+bt8EiatZhnPNV078U3fCD60jLk
fPBxsXYdVWsRrbdQl5HxiaiohkhYgHdVeOcYcH/HaOB6GJWLh9AA3mLAzIKeGDxN695YSheiSdkB
mmx6y6BMj2iK1w1i++7vJrGObq2vnjKbvEYqh2xBDQAs6F06om4o2Aozxrxum9JrWfLVfStnaZaU
7WxtTkbCJ8qaget5TTEd8nL09JFhSigQHDRsSHh0KNGR8N0wB8ZW2p5ofBp20PMtRvDKKxczl0io
EcyW1Qxv2mmqvyQllSNmpbxrNdW4Z1HzVDutz3vRQ2Fij/8F5wv8Zfd/91OBlbCFJobY0zPP+7EW
XXvYfVv4dFk2Qavcz3bJWs0k7qcpezRnpwLALfl1TAbEyz87qI2K6MMyo1bYur82mHfAIJlTfNTt
QiNaLFPM4DK25uGfIZQrJLZQfGeqYe9VZYeAWozQWycdkDF0L9Mxk4G7qBBGp8xBLqR/MAVL9aPS
/eAf9Y3DwmCGqBV7v/xwZds4mxRi4v1wVnvkyh0e1Oug3+KzYFTFOhiKEyQmc7i3PVvXuIlRatyq
7WEjMWuL6jEGn2LyBSB4bGenio5o8E1pvIPW+6By+JSkQxP/B0kTCdeVuuG9GF1UrJ+eCb2peFOM
2XPDREBvZ10J9OUBBsSXnYuYbfhiqUd3gxiYhprgNvVKz/I0V5G+P99ujKnzcnz4xG54ofov6cbc
lo2KYXT1Pjp/241ZirEGTCiN3d5SB0kvs6cqMtuZ8nAzD/lZPferI5F9VX6Sd8oney4oZt4QITzf
M3MCdseb6us2GCczHRNzPK0C/nKZ+Y1cKxBOs5C3KYO3lNUqaKOJzTMm0WttELe8sqcSjrlKhDga
9utpKZm1vdszyr/PxApF62H6+I2wnQNYc61tVc4rXDOugtJET25Me2u9CzBMfyMLxyWiC0boqNUB
qBqvPjCye0UHK3pK9+tpcGv/x5qxgZNdv+21hUo9ehlbjS7zkDZMli2I1WYW+Rfo0IkOZSI3nwdt
qnn3nGrtPw7E6ooJ6Q5wajjsURf8eZVeOz2uPLisWFqZIKI+pDSgIQoQI25VWK95b7I5aQ+3bwtN
Z7lT8nsV3tmiDvnEGn8V6nPW6XE3o7M0bdNEVGYf8YvflzQs4Xp+kBOvrnk00+oQDxu4haXpaFA/
N9lxj24iYeZpo7UIi2tTlFNCLMdb7K3JKxD76QxYqf5FCe04TJMwXKeDQqo/ZxxIOkkqjQ5qd2DN
/zvMAw5c+LMAM7se0Ei2IK92yeVLOkKmGqLWT4u0Jot6Y1nLeKs6fEGVGs8uepIltVv7wHk0SkLh
35QQtyknKV3b7IKINQiOCPfWQJaf1mGRsyuVGV5cdCtA3jpqAWLZBodE95djoKGhx2ioA+T8o7vh
awokx8a2dOw6E+MhRJIZgiUu44ydjJ/8IQ4FKIiCb3yESfPEMehlDcrBPGd73rym12RakmGq2wGh
bcwntaIKqkNgWooEGWI4oNQ+hHqkShBRIMQXqrNyTTt1wpEyBlk+W/clC48xZ/xXYnfBJWPwF+YE
WteDjdXFergebMhfZ0Eo1TDUBKHyyvI6+L8PWmmqEMysi8Vzr0EuNiI4rMnUulzsGWLfKfs+5jsQ
5dn6DA1knaJKbyOMsukHtyM7cINKy5XhkcAEGX51qbgttkI0ZS3p59TDpmmMCbjgZhYv5ycV7Cne
lqs/5DT+ZyxQNpijjemvMj3AEYLLOPtcw74WQdIbqRsS/wIsYp0MiZDvUPlWTZViQy6TGyEepaBf
CAsh0oL+bMcOXK8uivThn6M1qhbtUQyK7r72bcTggz2YnmhASoa+bbT5CgDrxcPbq7Nr40+LT03I
ripBcTjMnmoK+faB1o4Qw2SPaEgXENCyBuyZySiDdudpRahdS5CvqkcojXYep8QXW42nzSGPf68y
fYZ0efOwkXS1SlS3hU+SgeTjMU0y/qyFbznWjR48YHy0O0trHIN7mXIaRVaNTxWPyMpuN+eCiN7d
XPBLD6meIbd9De9Cci75CiOpqsFs++41KnY6wZeB0k0+LlHfOuoH6EYJF7Wu3+2CZCig7TypWdpj
+mjafmMxofVKtSnY3okPvQNb6zmzhSVkHc7gNc9WpM4zBEEMQi8WfZVCSB8dFzfRa0IgX7A4bHbL
rZDB9Afy7fJnSvc2fRcqCCuqqg2wNOG9nFM4Zgc9va4SSCjoRa+2t6cRPz9Pdt9VGWgrPfbZWn0v
aXpLFAdIFgrl/63WhJdw8PQmnubfK8c2HUia76piQzh0fveSfdgxu2Gfw7ZZqk2HJp5lSDq4+41H
MKBwllUaIkJkRnDKKuG1+odb5bNn5bxoJx0+Dv7fQcj//ZebYaXXTj5GVi8n0YAg4Wpv7XOBdHyY
sqqbz+u56Us8mYU07LG+XM2DTO/UHFcce4dzS242v6SNllD5XzD1ZEK83JHjbQQWTagS+1FPonWQ
VXnixSwt3DhM5DobqGas9n32eCQz5uF+e8WpFTvSh44K3p951ze2UfeiXw8VNLk6w8GFuSSG3Jzc
as+XzE2DQBhxG08uJ+lY5qE/d7SAJpiF+2HAdzWLuSttgilk9pwVCaaJUphcuYuGfNTXYsw5vmPP
FksXT8uGCIi7I47sRtiTF8Ze/ZoHKnjU7b8oOnHOVagP8KAGvlZvawqxGxRU1y08H9KVYaDjSfDC
gglTM3lOEisVZgbZ/1qPj+ixd5tKiZBcQj4/tYwsCEPPHfxrlBsOa45gF4ftuYLXiTI5OCpbndzl
xr5joChkwvRUql0TiehfSmqnweroq+H7o76DbukwMc6KOkRA8RmZuWIDc4ywdZAWAkS04WrqNUiJ
bPso2Ebe47OTQBTaWxS6+x/cA8/keOfLdbk/pU5ZF7nWXcqOpgQdsTs2Ejf3g3LdxsnpoCfdjgeX
9DbwlJomtqWov9d6cFQAfRwwFROGIyyDH3FbaC6c18AAKdQnmXV1Xz+GFHYMJQhBdCMfifezyX3s
v+2aOPLLa03ffPdTgUWKd/9mylNX8ygjwrxmu3DdsGLYsw16Rs5Q4tjadmd31voAXbsr5zwTS3H3
5OcRkVqd8yPhX6fmikokRVm/bJMhqbCqWrDdhbHo0gAZggaBuo5PC1WSTHcWusvP/+7MAOjQbdtx
xLO0ce5Y0WQWOra3PZYXuimUGvF5m+L2jyVer5y2vB7xSksrfcSI9GZXdRzSC2LB3oaBsWRclqVT
wGzCczo1carUFrN/APNbBdEtOo0H+RrCfaoVpVt8+aYoMKN/f/2wnSmI1jZwvr/Eh72EoH8b/iBk
zlGpE+dQzB6VCYoOw3f2O8hdxB7n2SzJYo8Po+yxEg6npr+Z8CiP/Cqtu1qbqGe768cF/xEfwNb9
TZVpfXZzDfVCfx+WjR8/VCoIWq0enK5uU6Di+eqpOjxYrGoN6Dmf5MoSuRRtgp1n4eNOvba1LWMr
xnrwih3nE25asIpZk1/AryMBhlMTctM4eyM7q4OIXEgH0Gkz7IwSTnGPpJoaXW2XB5l1eJRFyWT8
vdarPCLRMM5TFwQYyw3lQh5dnRF5QW7MQS1P0poT/pseXubZGGeCX6slOlDZ7Q8KTavzkUqwS1kt
P8pb8TCP608J2SmIxHVHWp/zZCmem0z14oFdSc/k4XZv1mE/Z2MBdZiSV/OA6wh6TaqJPAC3VQ3l
PY9vGobU+cOWddi9fRO4LypaJSmwjTqsFT7Wj69s6IQ9LiahlwHgmhvTEh9sjtF5ihnbpvovftOm
JlnyuwKz6u5gHKc5XnTGrFj4fOuWDRd1Gq/+UTCRO8+h4I7QD8Fxvx1VKPsEAWvPhLy6RO2m6Xvn
5bITkSK+brVskVXNOeoN3kaTI3issB7OFMRQ8RBEjl6cREXHvpDL57SoNE3dzckbmUENxUHddfK8
O8bzy/0bBYfKe5Ew7+gtT1nVCQMPGr5WTjA+cn6ec34U5vz8SRQtP4iEreYocGd1HmCht+g5ehHV
Ebw9/Zwoqs/P2R89X9oeQxVs/8178SAi+8kaYjY1bqndiUOfp9eB7AJgt+D8YDlUQHyh6094tmnH
ccgyiJT6vbDtfvml1eU1plY3QCGgyxt01uq2wcngx3mbTakpEVT848BSf34GxDTDBpjyoTSux66o
j8A6n1MIiSDoE0G6M8ZVfKIuoDd6xcjMAW903HAsl7sTxFDyN6j9jsDQwGzWfqTcmcq7qQozCplq
x/F4TU+d79fttrannwd0Yc3jdIDrUiVwQy2Q7V7HSFDYJ2KBYMFk7cFpCD9zitFDS5RqKSaGEOKg
K8E648Tg7KsL833WDKxZoLdddnS8ZhqtboS0dpE309xO7wE7PwTIAqd1fD2YN5pGuhWDQ0TsgO7R
VadZ/l8u55Wg7rmOFi/Vbc9l7uo2qb6zgwzR3nGHDBUR5pnmN77SqAxC2gkISoHPjaaGLrNWTDG5
G96WLSOoIJh6+K+3VdMEiI/WevawSNKh3x8F8nYEnYYK7ql2OuxcYqgnq2SIaNsXFYsMyhhL+0lt
NrB/xXbYBEPRis/guledHiv/sVe5d+Ng7y3K80F02PI21fN5roo+Tf+87l+cfn4lHZXdpCJ76QEN
Xt8RhwstPi/XEHxMtJHhvP3w9AM6oMZntz1KU6R0hLWzF9/eHLTdKETDGhqhyztRF98YWFGSe/Zo
LpKAOfmkyQ+ichaHZ/mBx+n8TaSLDN438yNdSeLmYjQ51e94SpQf5690O4W78tf03re7PIQ2ibno
JA/h0fqkS31nPmc7lYJNQ2z6MYTB/HTOMnuiV3nX39ukjf2ZIUhpgRlXIm1YJ2TV5M2qNEC8YSVE
sdm7/fqs73sOkTbY+IS+AQqe52sygcRR7Gjn4E/LQndO63EURv8eaUwo0xG4cAsDxppOdC0TJSQp
LwrPbdVkEszYRmkPnc6mNJ9W3xsxdqFmZpZdgfUQa3xxAkiRylLrn5XKF/ubXKkANekIf1sEMrCw
ioOkS7vvGKiTvflk3SL7GHu8FQy+MMfunhY/TTWwr3LKDBWWLzHjB+Xk1rnbfh/1qEv3PtsuqBQS
94RcAy3EXHCBJ/cYFOo3LPn4u00f6TIUF9G65TN3EkWEUEsIrrtBk18EHNmZCiQ47j1DudUVgJUu
ehu2EYYNXGnnlugMJABKIORPYMRjI6iUfeyBs0riNpatdnLMPuszcZDdPxAluAxnocYPxtHALYnJ
yGDOUr7die+qRneiAXFM8ZPtsVPguguMSV8bdi3UFse8AbR/FtAeiPD1Tvhkvkelkl2Wc2xzlkAB
+vGL+RUIDfnVYHX001E4r8RhvicVUoMCh2JlO37hOY6eQ7KNd4QdxUlqKBLTyhWVIoa8BvHrKQ16
TnSZqXYdqmtRzVuZz3Fa2CGDl9aYtOtymSXz4QBAqcDFLLz+WKZKyk0nrDicB53TLjDAK3dwsnTC
gmNQ1ytkkJJZnBf9AlZAviqP4BaP/hPDJJuB+WYBXMOnZA8JrXETCq3RssRKPgga/9yn4ij9nBDX
E0Z8gWsbcVxEMlsUgmrTM6sdmBu0ct/MG4jflHeMovHskU+NdYVnLOwTgJsDPPr9ibUdx4IXUnY/
vQKV1TQ41M1stliPs17SyWNU/moOwACc5I2E5m/J5757+NbSfpzr1FpTGMwJlGEGStREkGxP7Hmq
vrvBfHraedtSVNYd/zIUTYrZihhPUNN7/HLiaUBkkyjn26//W8952dUA9EKobob20row8ldkox/Y
zKPgA07qduky42miGw6625w+nhJCPjwUvLzliLN/DZTW2KwGXPzF+IS4OxnCDHzn6lcqEWgPnGwW
zaMBwUpITAMFatKA2G5LUroF8/LlaYV+IarAnPz0CCqYad2rU6D+TR8i4SbcvgoENXUB11YQwdCR
jY/l1go4fSE2cMrtRAek/sspnuDucPvu5tMRcfKhbEEFIwBVQAcmePedgS+Id0hp2x3q4x2F8X32
U6HUHymzeOvkCB/Il0KDHeVermkItWHZYd7HejDxp2R0kzVEznCTZSlmdZOIJNRK7YE9SI4BOoFM
UGrGUItp5VGDUkfLR/N/RkW+EncNfRR2L0xGYaTs82Y0DHXqH9FHOqzf/P+C0nfD0fttgvC9toN/
GfDWvFYQN34I7T+S//6BSl1POZRrVG5Qm/sSjQe0d4ZqARanEryIlWZG/AgXGC6oHvBZpj9wIOqg
XbDDV3h2swpkHs+E3gCHsKHURwHVBYQ4lMey0VKGWu97MPumfigo4SCkvE8d7YBQ6EqveaUC3la0
GtfafCR0qWdtVJkeVc/P12affg7LjLMBka+xMoSWrZkJYuvye5EXqZJ468javiPz7/UQbJlDxIJV
ii820O9gz4oMzh66oB5Pm6v6B6goAKiaIEAC7RWgOwbUp9ZBvr6KQnWWkDz02oAJHgAz45NWRlO/
iWrfNHdGI5lsuP7Vmlcj1SDxTxubHjyfNrIeytAaYfJwtvyFu0Y+9DyquhGAvawDGa7GmHKmjHIT
2ZMq4GLeniI/YhggcR+yBVPVdgAeOUXZwpF2c3Y2EFU5XeFPsKlPpsVvTx0JWxsLzws85eCS20Fw
Spdyz7ltk+UIom7xzyV5Ua31GYOR2dlscy96HF4gmNyZnlaPQHZSTSfqqyUh6QVHC91P5cfKUS1C
cPbMnmL060I8qZU6VK9gJDi6IiFTkNqO41m86gPQ9Ubf+c3pSnCAwwEDu+g3aHdGjm/DKmJPvnga
FLTq3oXPOf+00rlIcZsVqtPdtXiEO5He6WG6oCS79JNESV9wRRF7gKpd/Yv48QKZKGJLpn1h/Nea
UDnLBqWCGU0kQE/KVdCl/u3pXwf58jrpL4LcCbn2mRmca5iobMwjyGJDV0CpqVvgpNZvN56w5SUI
cYUSkg8hVCJGl/DLCFQBEt1KXwtRrRF/1UE5GHm/9na0hldSJYsLK6b/+3ZRXT/XuC/7HzznUh2P
ctVUdncSi8c4W8TYncs7meeKa2Kunr2zojrOirukhRexOY3HKgnbeyT3wYcA3gO0OgizHbwzy+yH
jeVSRO/r+KoZgJBiN+GwCUkNOMjjbx3+fTm1UjlACoFVTQy9U9uBCvIWo0e3m2ahiXNqTy9ebiu1
ojCFuJOcS4TX52zPfL1gZC1kBIluG5vt9VwE9GMgQiwITpWFWIIWvJ7qmxZOryscioev+209WVGi
IZQHfvl0D9YMzX+KOOJzBi3H2emsGp/mXINGviORYBz22ZviLzAmZ8g7MJLHnyxpQIUZPiisNEzG
Ibl9YxJcPMGC6aiEQGx89rVICED2sJK6UYaRfrPf01yLYhskzGD7+b9h+TlvceSqUePkqX8Bjel/
PxWAPwHLX6yt8pHBSvlCjF6l9jTxSRgCO2uCJbbVXY5lupHMGInDWwt2lZ78Q0gU1GuafkpY2K3U
UDii+EjVFWEqIasevuuDZJl4Lx9X7XmlL+ytakDhy8htvbg+pkAG0lZ3UOtv552z7QiO/wp4BKTt
7zqo3rE1pny8yppmC/kkctIeBIQqU9oKaMKPTHadseRkTZfE/VvjIQ0PSnqBCAP27zjkmDlX9XvS
1tSJuKfTuu2tW9DpwK/kUUh3ZfzHCigBQv/9IhVQXHT21svPP7sAMhVH2jMDRYGg+reAQ6kQ8Y8C
ZpvAAM++KJ4EGM5ETvNjond3WrOftfSC5Ge1+4r6TES4sFsepJgxUKo6We0Bzg2K0zp/DCiadAWg
LV4SBbvuPW4pzWqd7h8a6GiNGiP7lE+TdJI7UXqhDzgGN/nK5KJgO/ed1GB17spPbVDJemMwjUUi
jauB4z2Yft8ZRb8O5Oifdu8ix6gcvsEIJy9M+nNMU7OjZGfHpcQ5GZYdD2Xk6gvTeJN7QkYTD7gd
mlcVzbQkOdEVXUPTN7j4UNYpgTG74Qdk58uTe1skY+Mo63INuALWL7yAqXPt6IvMgFMCQtCXKasP
kzFQ86xrVehq7Gl3idtNDhH2BmqxfSDhY3rQ9XDVernqaketYGMppwCwD43HPgGCZcRIhnBcA4lp
Kj+55TTcwW7JxrnfnwLpnCsPPAxxj5jaHS3ChGAikADJeq4FYLvoxeQVDYI2rOhu5TGc4x9tKF+s
hq9QtsRsxpxE92N+GzWeWfmofIPjQRU7Kp/fzg5nfAyEOW5u7CH6Hd5nfFBW5d+fkXt4rYsmkXsg
6KkhQ70Nl8HwdGq5SoykBqmWY3UhTOfXtP8W0F99f/cK6TZpmceCiYzOFY1Adbk2SMKXjWEPAUee
8E9bG5ErLRe+raJt/HLw4K32Lk/LiSQOvHXQfKSrUweci1ae5LahgMrc91K0qwPla9FayQETzw+1
lGT41do8/1XBZEHSeA4PeNUuNomo+Gbe9VI/FCh2gWVoCaYRAGQxoKVnp+SPxp/VC2zp7JIMp+Zl
40Ed06hHdHmeNq9j0evjRIAT5iWzAQ6WOSxJIu/Cjct4fk/s9D7ddZR9Eg6EZMmmJjmF4A5VeG03
gg1DN6aj+XQpMqim7TR6hoRw1PI7nmPey44/PYaf26bC16IugRHCRHCudmTAYsGjgxPlBTj6RPKN
Jd363tgOMFjAVn+bAtOTe3bTKNoq6kWqa/Kcwo+6BW3c2c704zmmSXcWR+nGxOJU5THQb5pttY0Y
LF6UpOpieFrneiDtXB9pijH+mUmztL8AUrA+epwreLhmWo0eASYPh9Swi0T0CJhisv1G/W7yviM9
FZWdF0GQQ6j8ldCoZM+27zQ+RwhPlJpvMDDQKSdbwXzpqONZ/r4O5yQ/RLtIZsGHs54pV0P0trv5
KQl9bDOWUzKLGGNz3uI0Pl0kztI2M93scw0X+CglbF31pmE7xnfCUc180p1wwO7rQyNPeWHS8a4r
mRJRLbxnOlgosTj2/u7nxA87q+7z/KaXbnx9hqZnfI+b5hxhNuCu1g4XhhQ1uqfZYEfEeurFInPh
hOTyQX6pafvL+mg9094KevLx5/vZTN9Awp4vqwDZhns/SDo+loD0xAFnI71g2FeOCjIReoISNG+b
KmfU9vIbeLiUSZ9djEhhmh6gUxJp54evobqmjDgdQtyLZM0Bu4EZpSEEH3XpWzib6wLZosgUHJdA
B9OrYJEJT+tLKjLmh/ZneyOb980Pzwt7XaKRYL62jn0C2phSNXi0YMNcWUVY74h1Dyw3BbOvfMqj
eNeq+ZpjEhQMvkOPd3qy2/9r5Z12eripOlLk1VTLksodM1HFt2ZO5m2B9vcpgzSy1LFkRjQQmEtn
QLyPiQnzkyblsu18RQXtki+4cYKfGFytsPS8P3ir361xnxuLZvkMwbqzHI2sqhRRd4bDHreas6U+
UKK8kClMbA8Gbt+wacweVC7pWCg+AHLLeN4RLObGSMeRjDmi9/kNzam9piINBTquM4kMwNyA6wul
2Z2N8Q/2xFyYse9HJ/Gt/MiWJ65T9/OZETwzku1zrmT9Rb8pMtaG1FSdxD0rB1Bv6JDNYCGchkmZ
3ukPuPK+hfoG9A2m5dy4DrGQh8Bl8L+VGBQGmaWA4T5nxZ7kE4J/dEjtOGYr7i0mgvJvqvO0g8az
BOIDf8wRTb5lBJvdC2zsvh8kUZFBdY6qweIAT2toSyAb1jqJITYju61RPTIz2/Q9G/qsw2iiRy2i
qalgzMVCw+v+G+6kHJOqZGNFJwwu24dybpjk2QR/OXZdG6l1tHhuiVif1AAJ2PQBX3SJSJBvL//S
lZrpI0WymOcNOdV3TJ4SZi9d6BxWMg/lcA5Rs4HiJ5Q9dQA46v8BhsSyFsLYAzNBAgZT+RzFnIWf
VoA+MWoboOHyQWOMEKUhbpbJG52wvAPl3TbnwxzjpRwa6fwtC+541RJP49VDJSDWi5q0DzagaMyM
rGD0lxj84z5aUdrzEf+pjQ3hp5mS2ZEcNx4i/Uri+oJmDO9By03NcfpxJ2fudqZUZOmanxaE6Jah
rtkA94K2mrLw6hC4gxINsM8xO28TWSqxtfzDSI2zt9COGHSAe9cRleQ70/YQK1EWE1MKwMCKPry3
MqQ0mqpp420CkYG4tp0Kagt1ArhtSklSb77XGfswpQJFrqgnhB8FFJ28Ids8cJaU/CERc1zRJgap
M8nLx7aBuN5poBBg2epZo/a3AEmxnB1bny1CleV//SQVH3QSca27bMVeknYTXXAh0pHpCtW3ubBi
25nXMkc81caVHcglsTq/Arjyw5R9m+9gA7Cn7WdxWsTn4MNMuWttK3ehjzrYutHl8DVywa86p0gN
X1yorOoRKipCPWoawoNg3jVqgBzYCgWh2JUDYmitQXJe8R7dYgWBvC5IKYp+I55G5f7uYzsxQkCP
xntwKzanTLo1TPCb8O7I5p6jP5TpDRHNRSXJyaShEPvo++dzfKQKHJMKFR9DRDk9trzEzA9JUBcb
4ZhiBzve42IQ9T2GMHY1oJ936wEocAGB1NWTapvTfz11F7sLWya3sg17TaTiHi3IcmSzZXOaNTSA
xOvIdX6vIDvbCXfVqrns3X/rYf8YhUJy9Y4C6xlkh94iIbfP2/sBfJk3nrV3Fe8OBx5MV57WvS04
+YEkjQSADJDrO9hemT/H7H2awFT366WWAbcmI73imfVP38MbmCou7FkSjioOvmC5U2zu8+3h9bRv
E2p70Hx0IddhKVxSkUGdjm9r4/Fi1eiVWiihTh8keVNfleZS+Yt/YYSzJzUuGZT/PSCU4N60LGxC
noXktTHRifPl9apaHQYNKpJisj6z9MA+LfYUcxmfY/Vknw0kssPmwcPhgSi0hdq14XpugYdOZhT/
k1kQEmwJ3UDLGkUdqnISWgqsMrN5X3yGvBhI/Dfad9RUBSZutwVmuUjBwfCqeJMD0GVvxk1bSD48
zq08iP+9qPcf8r/we3OL6tdfsXMIgOsKI2qaPc3d2Ea4PDlslibJ7f80XZe6rPNIxU1NcYJVuI5y
HXPek7WyHLVCigvWG2VLs8VMZU10A6DxEp5OaKY7c1NwQuzlqoSIpXJy3f6xdS9lu4XSoLo4nuXd
hYwSSno6+d77qpnUqpH2qjWWzXpY+tGwyrmKqeoPd004rpLwoCU2V2XDmjVSxVNcLtDSH/TLCnsc
2labLrSZiZ8YBBYD2xBevfjgKXZMJ6ZKtabWtvQGH++lTWak9RAduA17X7w5chSLBP+HbwMhDwNv
v7cNqBEA6iRZa+tU/j0vPDfLpokkTnjerpB/lfWYnXOQy7A/U6oocktTbx7jIZ5AwHfEIpGQXcyr
cXbpyybadJ1ToiMO/AohDUXMmIdn+haPrOJpfZonF12KuSJ900OKBIrFtGxAaGhxgle9hNrUdJ8n
ZAlqjEjOjl7cV0bx9wLeV3ighCj3ylyVJkCto/JpBVttKF+PEr/VI+zK0BUuqVjQqjOHAZlL530R
91zNCtW5lZJJtFamW5JLbl06R6WcDEYUMufU5OXtWL4S/Dq6gR4r720ham9bflM+QPsKDXWj7KNp
0b4I6/1ukERDi90P3fXPX7hFLIJBh8QYlL/XvEM0Q9YFSk+ORzhzGZYxbwjUjmjmkfo5mWMqvkNn
RYR+9alzWqCQ2YwtWPwfdpzfeEN8pbR5W5c2zg2DYfSBhTeGopCIs7JOw7YkU2RmjO/aqjlAR9B9
1jJlFt+N9RosIm8o06TSFNWYXjBBdCsndq5hrCIdIDeZdbtabVjCDM9dOVBSv32Ag82NnEkF7NvF
JkZqqN7k0RpLoQ8Pf18rRXtq3FLCT8sl+wdKKOmtasuREiHHCvYStlrjvSgxiKY64wst2zYWQCl4
9vKxjmoYcc5Rc+xfg4BCzhYvMGmADgPUyDQFT94/O52Vh1QJCsOGCoU6Uby8LgSW/Q4kCy1zDnH3
j9ErC35wxssGTDhYDxyj67epRQi5ZLXoXEkPEBcRtXtDhphWjzV+VhiqJmLzba+WIU+RMYx8wDHA
Z5CTd02+gVXroxcMFEfLcccGMynLg1aD1UVSUASTZEv68pbOh0v2rcqLlaaPOA2+px9X5w+aGxfu
PcP0+QRcmeJLJ7FbFI7LXPBCYeW3MRML1QrI5n5yI9r6vrgQj/lXtXroOESXLOhWpb/L0XZ6KRQ3
coyravIE6IfqE4xYlAAcjy5JhCyFFnW1dOA6bLUotRK8jk6bTk9pHxmzLXC5UD8cfHqcwLwRAGu2
n5KDgDXDsDEPpp3skD/pwuvQ8VL66REyZF0fFYC3CY4GHbsf9Wp1W9DAiOr215LPFxf+kNcuhGIo
mfXzPMYN+yqGJDYSZ4AoD7DVw8grGElS/ZmTXBt9M6HyAWZApPc9cm/+lqye6UXpfQk4at/1AOsZ
TqjSwC/iLB2otHy5bWVvJk723Vuw9Mz6NGYoJI8vAtJHKlQu0XyF1I2IH/0KxF+Bthc1iOHYtW8o
3u/NepGqwVaKkiYZppiKpvz0/uW/hQu95mPQqpexnBPZBX6XlZHlu5p19jH6ZZn4h8Zz/sIsAfU6
ivEwXvnLUnus+LrVmfpUwivrtPGyBuJTkB6bGfaQvbwitiHeb24DZ6o0FnaEgAImhMxTUvppqLOl
xrSwiT4+eTAsrS8WLyBSbXxMU6nNAEDm4xVqpr6/AoiPPO+cM5w4D9iHcGPwb5W3MBNPQbEXadTX
bGp/F2fLrN9LINL060NyHKgpxTb07b7k58WGFIL5oyNHwSaHrTR6n1AcTvCy3Lu1MvMmzKVhjQqW
fA95smI3KNYyD2cZQZX5OJN3lPV7FoykffLTLJ4Nvul5aDjMfe8fkS6DNWtDBt1Pa2aHHVIZU5ZO
hLlFRh6JgdrxVkoZBY2+8Y89YN5r7+01yV17qkgXnXmbkvfsr3w4KVbREKkWxjTtqASfjlU6g0j+
zwkKKOSUYbCR2OXr4l9ceO+0ge4udP+9Qzb3stBB/UPD1suakP3FgiawwMiAC2jW/G2kiuRz9Zup
BbhfV/lDAWuGw09GR7MB9NEvmD9hzTaABii+CYnEkjUIJYEtge380EWPR5U4r7dt59t9EDr9h7WX
d+gysGv3B8basftLAWLqkonk1RdY95uTpuSZhxl5KQcN9zS5MyUte1ZRJPN7FPQVn0d2J2yJGh9b
oE2X+gQfNUhme/LjPyXvSlCscB77okKwi+wpR1RSpI1do+Syvvd7+ejwXVcPsf0AOzugs6qwsRVH
myUriWsfF23aIuLGEX2Wai3F6nw4+Bvn4Gj1Ym4TOFiBzwBWot901+xUmilUgutjDbL25zBQ+TH5
bZ1hzG08fb4Og/wrocBIEO9qBlbyHYp9TFY9wKbqAMC4cjMGDUOozT6Au5SkVfuANcGqTMzxcBFA
hTXwSUZ+QVwM3bgk3ngd4HcnMzQS3FOh1eGj2pMJfIVkgdgwPUyddLGlAsf/CMLA/yAYeG7SjWxg
aBVjjoarbxQTOU81SpcnIgi4A/ZXK3N03B/LLTi15oTtNRCsnRsPBwXbKYOMsGYzSPClrRmEHHK+
nutW1HUNBYQMmd0KZSHOS4ng3UYJ7bPQ1BhQmupfyz1IklQZlW00kDivq3J7hL1EvTDq7/nj6Qt9
1988B/+hjvp9eOvyqnn1BqCwEwqwE5AbAoA34yjBhrGqqOf5ddM/EvpY6lz4oic9J9za1oIM5Wzu
SoEWGYwYfsaD8k0seyhngZD0F4MisuhVvLEN2BFgsAnjoUnHWJik5DAlGjVl48RxKPKKb/f3CIHc
JsXZYVftJsj0V+AbGft8SYdNx/w8A1ctnEZt1Hs2EHz89oTA+TP4kC/TY0vnLhWwYsNCy1Qffxjg
QZvJMwC1gxwGtldZZWXX1NFbvcXfas23Il4FJRCDjzZnfuccuCJe0MobMvjWOgQn9gjvay9Loooi
FbLX6Di5KnBNo1lvynMiJrRvNT03rsRr3D1Vf2HKVeCz8LYMqSzfMM2KvvBulIjJC6pXlKRZ2Iyi
NpKydUMTD1mtKFosG9KURMfdvI8B7qbb6bZiC174gxS0sz6tfWXL5yLv0PwVXuSyGOUIG4GXXwYc
2chzoW2LuLn0tN+L9Ti9OOC6aQYlAd2a/WLVSqYQvX7Tm3Qtt/GDLuhdpIH1l87FKwdYIuQbl0OK
kSY90I+XPTuvHTCRjoG3FRCuWtCtvZkn9HivgGYKcJ1b9BjJfR5nvCWu6+0q40BQLC0PrD/Q1wRz
F4SDccnUjWIEYdp4Dl7MZIfXXsIxJdSlBaBEvN/TWKS0r4keJtgmHVcHj2Y6pb7ApQYb9hA/ljWd
xffb1R8lV9+3Bu2LQMJNU0qNAmM7Mzvt5CXOG7sI9p93/K6ujnkoRl0mWQK2G4mjU5RCIZUtpimY
KIxL6g8hqSLdu+VuWFoP8lpxBXwA7yzL82IM1mTtv8LtABew/W9kECEMly2zZIr8Zb1WBMMa9zNP
WCo66XZJwyLmeHVsr3Ye5rbDB8cg0I2oPvMm3665P6lrieb+0x6dckaXn91MqWuRm4VYNxAOJpv7
aWZPH3mu+0fMwkePPlTjdRei9SZsv1eRy5g3FCDCBzh50t2v3lxAQXgm/WucunUO30NFkzaIydfX
TZlz20HVkM9ywlXkaGC0gHTIfCoiVS6zYND9fgno6rJSVKzbifgINcBSvJdGstRjQXnJ7oeaIR/F
bv0l64XbHugh0izvd0PwpGDoDX17hZLFEVUTe99Ri52NSnkhYaHZNsRQxPCHUelINXkjFLSu9Up9
j4ZXDOM+YV+NaOwgA+jjdHIGx9stbptrI1ROiWUm20jryZebiIrTnoz+WyUnW0LHsyQYMdq71sxT
ggHJvZgI6OYhLmxqmKAB82DWEioNqJsTntPtqAJcpTWg5158xGPt4/VtURu/uo/tYK7Z9gcV0rr9
8lORVZG/7Bmvf24cHfTjbna5sS5ILNNJJtB0A3XIY0vO2lMa1UXhVfCSsQkM4oa/LVFq+nvjbWmM
iq/7LnMKXTmWnXVhYobAqGaMZrjZ0WY/hipTWWH2gxM3HfYKR3DZMTxToqihPeG3D2d3pP2YrtJq
kOB85eJNTItP5DiXoEkicbHmPaFvO2XdD3Gw3+LnoJmbqdxoKbeN9MlfNfqkAmh4yFEZeoulOVqa
MkJWHlTC+YYanksJIM8yYL14Y4D7lJxqhff81HjD0ieEq2yP5TWB1kqc3mg32n8YK0APQHEuhX2b
1ZyxnbPY8sjbLezcAtj5ScLsn8BCCZTEe+yKAOfDIL4P6NMbrPpXtCxfd9dBeFkPmnsLPVWT5kEx
L89EeFAyn3tn8usKxPk5HUTIemRejJP8SA9TFbxwnE05+fDLa6Oa6/f6dcKjI+rELBCMmAJe6tSz
xfV5YEs1NXQ90eORvX6FKupsTh4b5Eei08Di+eZji9T2WAeHDCgadbrQKOaryXwYfpvwqz0zVIag
b6BviCQXGAsdBewSeTd3DkdecBRBweL52pThbE4xMuo6YsCLFRuGYCT8gEE91qwYmOUBq1MU2CH2
tv522vdBpPw1qI1bpP51t+4FrGEq0Cg1Q8G8vfyfy39zFQs0EdEtaHlEuiQW0XEURblwLYuoLIIU
ohNYZpoopAJixiu1ZOeFPKJkssSnMA3n/RdEU2hL0dtLEwbZiRrI8eRorANPxxvFLRwbsowOlVs+
aUqEHxyRyief6WHXOMBn5X8uuP0KuWKc+PhR6ViZr3G0tfkg7AfJhsKh3yg2tUEj/MXR9soo0+wk
BOIQoStW7a0uAnLRm+LU5njne1kNpK1lxffjTpFYuI/ZtlVOa0X1X5l9bOIvbF/0m6/LKkxYG4OY
frw5Liz+5Ko95lGayG1t+RBnTUWlI7hv0DVUDU5ZyU+dFN8Pj2VXNBWeGtjiA4Y3jwcG8lAYDwyP
9gaDXkGMA2Gzo3ggz6d37Xaj8TvhBow66hWW22Mi7rALZ7TfEv0i8Y+N9D1czG6zWKIM40XmSMxC
5MP3EOxM5qU70jTgKSNVM7EQh7rTslXu9pBnmTix0ZpwcqoE0dmpJ1bVmkR7faJScIAjg322Q8nb
PqfWOV8468qRIDQpaH6HXTPr1JWH8ZsJ4/FNgaZ+860VhadpxmW7YAgnQw9PPZ+1vtoWdfx+GF0B
cIFUl5M91hXeOZ6UlP/Kt462d3nkPzYJWtQLXeGPEYKycMVdK9gbw7KkoKX45Fd787y0WKlZ93JY
yT5C8OkMZSTsVKB2bAL9Y8kF0McCKBEpLdnVh9y8HdeSbhUYYR1l6KKMMmLlAkkWikTIyVxpAZ6D
eG072k5urUUstX7ObC9xGxcqXe7g/bNwNwrhQY4B+qczyenNO+ZA5+nYkL9RQ30iT4ma4cW4aBN6
jbPbcqccMKFuOy8YiKvbKKfIflohhtgCz+TFneCK8/NIbmClHWEyYI1vjlOfuVXv92mt8wInAgoA
LzhSsrTIhcmJb0zDbyjYmTykP5cdv+O51H7gBe2HqaswyczCqX+SeODlKfkLMVN17byLgs2Ku4C6
tQ/uXFvhrNb0H6crfaxhC5WUE1Vg0GLZq/IIN85C/XrgU4nUvOT70CCaWKaarwMLjfJStRPJg9RN
FGCPf9toexeyuw2R8U+EsD/txRziet/CzTZS6C06gPI7QAGuazhblxwtDegTs9nLqOfWGwLQQvJE
mb4JNhi5YZSN8tcIdyEAfdpbI80JIcChQU7JFSL+i9daA++pKhgD15RIg1jhdBAHwShRJs4CwNi7
qc0RRtvf4BbBmfiC74x6yCNNYW7VYY6d6dl3jUuU5RUlQZs1v7KDkyp5/u6r2P1XZtd/13qGwCqT
T1UsJ3/xrrbo5U9Kmiflk/OlR09kD/5LT7EaYMAKOOBLpV0acnt2mYLbih4H4wBCDfaoSd0SXXaA
6EoiGG5JwU1ANLWDnn4bfPzxf/A5CQZW6YNL5nLJ8TLBsUAg6JdfUjVkn3Gf4Pm3a42CxuWSLVEj
AcRgzSwa2lk7WfwN2WCGWLVWUguQUvH8m1Ix/klpXaaIeeLEo6U6QNRQFIk4oMKSoyiNwjQca3im
5ixPbdZR0sRr460Q4ypQnFEJgFR8b6tBvOLrMpxr13tliK26Vx3a1/7vMv68wMN/iCDL/BSFh08Y
mENhZjRSNZ7/hb3OrL4retBWtweV2eKKhaGvqTyu28X5uYbWRn88uQHtxr3+3mV4dHHl51BGvQbr
i0gGEIngy9fPaGig4P9SV4xoseVTLKJ40n6SXvB7/iNt0DIYa5x6fLauSVdk6zlZpEbpygCOyOPo
zwPNBdXBNo0k3aigRGtaej2yCAW9YouFEvGgVBad2DzA+09ZI7tAkjINMMoSL3m7qwkci/FQn9wE
ZLd+DtoERBWgZo7kypSPiDdnj25fxD2Eq5SvtFVJeZSDw9Nq8UWC3lTgKxR9BvHzWNsbZjR2Xfyt
VNTfO5ITK3LqlK1uLwCdP3HsbAEJuhsP4RKBi2qr+8YrUYJNWWADSVXjcMAm7IgxPnVIP63z5bPa
lrRXpEbuHGzJsUdYZGsUF5d7my0vA4sE3XN+c9IR20FE8zgRDyo9wDeByAET98PVAVo8Rs+IphIS
8kUA65woxecP+vyn3ZS+sis1H7KqcLyQnkZPAjoOTD/8zyiVUt3XXejR2DLsh25OuT9E1J4g1StL
ykWrQuAb2tk2miUchIzqzqCOy5htdx9H9mNzDsxDZlxN3AMsDX+aurX1G+Hyx3liVmE8r4CBZt0w
th3wQCs2Sk3iJzjIhB4jzywMuydmF8SeLsyoS0xzqTXpegJArrnRmpfW3mMviNBjyWphwLuZBJyk
YL1PGyzzrM9n91zZUIRwhY4AdRbd2XuN2tMXa1Fp13liGWk2SQK3pRt/ov7oIycCU4lVUwP+4S7o
bhgAvPGiyDRXYWOf3/HsjvFHivToqVy8uUxn5zYqGLK/cFATWLhgDRbemcFcVGj7BRoOJx0DfEDO
p8bjgm0BcZk+bplTRJJA3jUuI8sIysAji/LKZri+A81fb1MlV7K//jvCfEpre4i8YQhR6ylffmZD
KN0u34Zl/o67Vyu3CRzMThWkzwkH0Lb3aI15WwXiRCEL9ojLgHFJ4ts/lAUSQhTPfXSFZer60IfI
VXqEzBLApwXjB5byAQZj63pUdH86yBIvUfQCToJjp/dL++T98jvZ7uN7I8DRVxXLm7ruDTJfSUv0
Kx/HLH6wFXAUNOpMXJ/0TTLlgJpDvOgmW2cqtJXizLObzpdxcwICIyB5UMwnNMUxClRIDt1/QdpK
RlWexe9fwF0AViE8y8eTuBcLvSi2e6YHXNVn8OpFl7pyNYFm6bXsowOyR9cLxizUVezDtOPCJPbL
7u5G8GPdZnE/sZenwMUDDLZJy9rcCz93VJGzsI80Yo9Kzf45ddFW6PsxnfCoP30fF65kG6/F4MSe
4bRpDaV9IMEkV6kV6qFCUz3IaLPYHKmuLBG6VlpiOg/s1natzE9ixj/WIx/CoZEq8fDIA/a4yEN6
dFdIEXHGbSRbK6gfKcSS1v9DNXTm5OFmrcSvg1A933XjHL/HhqrMIULomJIWWCtViDoQhN0hVo3G
j0xgBTn0K9IgK52offzZVapyB5EjN50XMYbRDXrcMzK4fF7oogki7rY27oDwZ306xP/xcyaYWQ9c
PooxiH8BpdyEcTAXOUSkXd6CJfD4L20D13MDqxYbaBZZn5pbpH8UhaG38Q00l1PTBCN3kUc6tkud
6r/FQKH5qBhE8S09idWhk86oSXpbmtTK8o2goKnnxY861ayz4fj4JFCNDIP6Cr1Bxf//J47ZYE4B
1kvhi1MDo0gkhTff5mRAFg4AZPOVz1Xv37yMky+HnqVUbqJBPG6+LhuPVBsIOJWYa7Cqizjdrx/f
UY9fmTJysai7tv6Z5pCJ6Hxb4YyECxGXEm60pdud3mkTaxBcBEQiYeX/Uol7/XP3S+UspiaXj+D+
rxKOFAMqA+PJQ3vs6jJCOVWc9wBYBWco3se4K4s3fDd/t0LUhBJuctinvlmhwK4HglJCFyfKx9Am
pyV9OFrIrZggdEhEZaDPkOeTJS4xuWNrYImcx4e0XRXuNTcWa5cRRr+OuL+8stK2brhMED4zO+U0
N1odPcnDdbnOg6hhb0sUFVURRCAc+l+CEkAOd4s5UyW46qXOY77bkMrxY9wAbZ8bfTOp+8NdeE4H
cx6LldktRdbH5iCKAQ1C2rPiYpv006CFKPXLiXMY/RdeBA5HiZrqPBmaa+grf7HPEWpKfM5xZXsU
1mH/nBup7LQ16jaaW4SPYXeU2bskk8xufpJA3+aEkZ1C0c2m+jfFJqpvxboXGMF/SRHid0Cqr6Gp
/tYfCM/KGhz3WoaRGoQA/vImI74lS38B1j+sV95XfrieM0BmDFiLrM6ozzQecHLo3lFAi9l6ItiA
DaLUXBnSaHZzee5dDaDJ/7e7FEa4NZGI6jgPdev1Gb1dclQdgTxDo8tLhCWT+nBbrNRSKm08zOE0
iAizVxn7Wi0gGPQVcHSGuWHDpjlIpx9Ld03z/mdGQFubYM4T6Ua6XYcRYWsYNsrlsHkkpfMsFlQ3
lh0OAYoBMxSuvnnDhwKrScFtJDg1JNKef99tSceVy7XftO8HpuwkJr9bM6dc90keYES/1Ekk6TSP
a0wlUDjGyQRotFP/oieHkc0EXsIsozkrTL/epc5xd2I1DXGpHQgvTNLqEmAZUi0+EqCjxQL7KVLX
1xdlpuKCMJTwO35WE5d/Ne7hqQfv7Lm+rXqxD8kCjWOWgBuHWbxwm0CrQP2JDvhk0D90IqQFNWnh
L5dDq5sp6PQpBV2ys4f7YPf9qZNttWt1aTN4cL5khWYXvXs6dN8cWGb+9mGXiykeCrQXTM10y+WD
DvCPWbFYV2bpEeP7URkN7lkaYJwYG6O9EFD3Jgm9bMztkQ8lIrcsbw60YPf6vKULuT/ko3ej8Gju
pBkKOCS1YEIANpMeyzUgkaS0wSXe6uJIdPzFGFKwXMsK1Weg10w6yhJeaPztuOJXGWj/6zImHFN8
DABp011eUGoNi7UiX+OZKn0zfUxknOwfVaTOCVS52y7DfJP71SxTiGvhkEE4Xv+3qvkEnPKFN+PR
JmSD0G1HI3iyqlVpksdO3MXneZD88Kgx4lETyozFzByHrYe7EDZSVFuwn2rcWBUuSCOkF97DpFwq
vLIZuWvNi5CahVpDq8orRCuq4ZR/I59/N/be5Kujj7x93P1B+z/dHbupx+ZIL6m2yy+H6vPBJ6eW
qeIjoHX2VmaGgp0FTu90joPyDwXpM6wEyyXf+iDlmr3eMq/GFCDe6ztTrCVgcRt5dcCJUDPVJYZh
vhqz51LJBjjC4WC6Yp+rrOVm1YJxMLghVlnt/XeDxy7XJyH22p0xH4D8+e445/l08h5BkzRJYtgu
y8v9nJ8aCOWe9odsNkrlwY7do23fUP4bFQ14OIAn8aoJYu45a+BDwIfJ2N2Odqj/w0GNblwG/Ii3
m85c3uWfjIuI4XLUwWCdRxP4Y/sIqX/Ocb/jaW6DqtmzneRcyOaBHUO+7ZNFEowxZ9qfW4EBScMU
QWoTJoGt5civ5R9ZgAqyS076nckVMLrXUpSdzJo/l/lm9wsbYmZ6icG9BCEa6y+SrZbc7QwlY25h
+SUSZ3XNqoTw3FITO0bvdDWhtvf+/NucB3ADYx9BhNlFisYA48Jl0iUtUA7Ktgn3yY8rEXQiI/jY
YEZ5+gwhVkLG+71v4WLM63uyvhwS3k8bCPhgVIlhUGS4we5xSv9Mia1YiUjF19E38X55/0sM1ykp
LIwK8CMsoh0eexy/mwZUdq9LYkMviibs23A8TzWFaFXMbZS8mp4kIG58/KXjMGrOdG2i5mmTyrOA
aepvKPjnAW3SyQrlJ0WAGFoO7MGAnJZt+5LPVVtmOo0n/KjxA5nvNybyrcMuxs9ojmYzFj+YI3Ad
6aAujgHenKv1s99dL7GEwO/BfNTZ2j9ZY0WqqQggKTt9jLkANHyT9xDdOZFZcwx7hiAJ6mLXcGAL
21iSY7x1w1Ov+ua2zcXtIDhjS6KlH4BDZ0xgfNDD7VytHpdm6vKSUyXO11AU3AB1VekZ+kdrRp1x
ZMcx9PqZXeeO22Gvp3FTMJ9FZ5fWGE2/rQGm3FJ9hDU8SHj+r13P3RZ5IEXoPIuCrjJhMADGyx3x
AAUxJW54U2qwxflWqUgSReuBHSYcHf5MmYPxQWu0kjm/1I7NzcY7kUhFecvPbeuofSDZb+INKlyA
DnXkWRZAUFi73pOC7nV5xt7ogG3+Jxqe85EC52TPmrIPlYSO3ziTjOD/Wy7ny1XASuDUOxKQbA53
wTutFWyZiBNTmTNNGs1UFc2/BsFBKIMh+tiIsacAh/QxJXsIOrrmhz38YHj5cKqYrwXUACyug+iL
YoCdShExYB5HCAjD3OOIXGM0f+ZtbFjG7pGz0m47PAekNu625aO2n9k8dsPBb6ILmXABD8/S1Av+
XHJVgU585HL2Zy3uWzVowY9Jl8+Fh1BTO1i3arUpH1a6xM0fD8I4nMRQt1h0YWFpWbvOChOGkl54
P/9fC4hVNbW0ClqQ3F449ssjKEJql8zqnmafkXWcx7/Kil1IQQfP0XEgQ4Bgnnw3nxVyNy/IE3eM
P7xoatdj7FwdmrYHoaUQfYZL2dek68wyg5sYCx9FME6B4J47Wz84i504RuJ3UspP6OQ0G8RKsNC0
mhwGdvU0Dy/u5+BJKTmwqM/zu9APruhpL/QzBHdvACuGt7tvpBkKyMS6+uTCfVlyR/Ym2La4fsO7
7cRdmVRdrHytM2jp71DQ/x+oFfo5PTl97kkMJviD8sRW/luOd678/paw/XW03jknYu3QrCQ056BJ
NmW8e7XfNv/dccdGhLxmUPE6ZXUIwr2iWJfy9NsAc3UuOG5dqcixKocPCJ2xYOaFn0MninRCj9Kq
fAH6CmPyicCCjD/ZNQJwJnL2C3NJJAwVH4Q2tG5X9Qqp/1SS/un5f7Ru21qqZ8OeYWUIakREUAgP
4CZ+O9+3KI/5c1FfFYA1MNWmQY4rtTJIs3JKsRM4aGex3QeUDUI6f8R4yTcj/yp5yAku6IfyzqNr
6RU4YlOcsU4mIsBcSuEGn1wIfCovmWAnHyoX/2Fe3PYYDEBJV1h7X8LI79x6RUkxuPxuf5DhWy3+
pLop9T5AQMrQjpKjhAgRSgj61cr2ELv7oDsy5VxlMtNhrq2Me4zXolfpPhr4PzdisMAWE11pNV9m
Myil8V17dfB1vIUNHSAt+oWVR3PLSRsKgRaoGmtKCZSrsYQp6cyoqxbcNsjdb7S5v2XXWw1aqSfm
x0qB35EFW6j9O6gbJZB+Hevk7Vpo6mv/QeDayvRp6ZdAz4im05rh5Nb3pTi6pOF16/L0KRHMIk+q
woYU/nerp4BsdUrcC2ApK8H7b1dX2R3KAzbFMaATgAzs0GKesDEZjjLP9Y307Vygyb5TCLDu/9T4
HVhKNY3T/SJnVBMiOTNm8pBzBNY9+ZEEmuVbbOi9sg29j7A19PDz8qCJjyzHX+rv7gyDrb+nqGNM
f94DljfYvENCh3ASMkTk/57qiJtANBTp/5N5LRwesmkrsmZoXD6EsCDM2HmvqWphU0UMM2OXoyOF
FUZcX5iASIRGZ2Q3NiTkXa30o+GKyju//2gInNrfjxbEzEPKAW88A4Hw/kEVaszkkdqtNtwOn6YK
0hXAk4b8lNZHflQ2TVYemq9rFHD29Byjf2zf7Qx47U4HHe3KUBcUuuh/dG58JYNWLoJ9DWTBsUIL
6QihbZQxGAd5pjRMHOQ59ZmNvWJyKwctWarD4lJYhTlaVEAxYi3FhuZzuZj5NTDmErlebdn8U16h
Zo0whTKl3nvbWMacq20h5OnwekXCWkbjSqhYsO5sxgvWzVaWMwn7+seXoT114luw7e1OoDLF3RPq
GWjJqgtM4FnFBrrvxRMVKoQR4qrHsRkINR66iaMH7/g6ptpg7kPlEyWXhGg6gL0KFqaKujrUgG1h
fomW5IYMABwMXU4gDH0ncSbDG3PG1ipWhuq1tkWcdxrjYt+oSvoobGQx+FfKOdYbqJDLX7zwy8OL
0xfF2pbWGEHzhQ1+TDCR5JElgOvKw2jxrM+BceRbqHeLI7wvTiOefXX38bFzq3/JjDvgsRqTqzhe
STCuelsiZKuM/T3nMSs4gqk6q9Tj2l5ey1efBaxG0kNhL/lMc1Vc2LK2UIZEKahY9KZuokOpAS/0
aXTpWLm4z6tRxw5gKwwoCUZygevCvMHR0+E1MA1MB3gy5RZRFw8WJtS/BuxN9eI6crsCUeeVmKPS
4G+90Vq4HE1vp+A/HejwaejN30ZfzA43d4ihmIjNKhm5c0O1+Spq/3ZBbioXweoX4/hh+g2DKPIV
pSGPfXDfXoDneM96W1+Z0aWku/BTTfbgQHsG3DlHNOQ3GVaous+2NNaoz2iJKvkioMSqLjYk2XRJ
2anRnDip42sdkZgueTThSrvFR7ZBDxV0g6w10kjpi5ZMV4Lx7xr+IBpMig8e5aIJe1JNMcVVvzRW
okeUcauHNltU3Rdq0tMbIbUV/vvWiQ8k2nZ/YcKLXA18JZ5veBiGwqTb8v5eVfAQvEsggl+tFw9U
YcIKtdopBoVLcTANnJv2GdvOw8eLRdCJwSvJqOtf6WNaQyNVG77cAfJ4KGO8dDEd+OiXsa9j+VED
mp5se+l9po/WzUaY/8LtBGXj1qUbkM9pNqHQBiEZatBGjnYPdLxhhGeNEf4tPesurYxTBCdRJOUg
qbxFC11jTBQAILip5HwjV/JaCLEqGoBYEPASxPNBiS3mzmRm6+pdDZieqI/wfGhTyaO1R3wE0ex1
1pOzqm/L1Bph56hRwSGn9c4CU8L2WXTgJ+TeJUqv+KECTFJs+brlb+5VPI1VNxn8ApZ1ngZGiMDt
3HfCvMa7wQ2mr2EUJUVck7f7Oj7jSrEzTGOBdQTR0LHOOl6xe4zkCKvIU4IpK2uPJ53nW4Rkh1Pv
9FeVSA6s7eOYgSqyXUSEIsP4KCjYgN5bg+0T/wIiXGaTU9VNt0aIi3p1KJ5wsIlzuxOCKaMPsd/v
XcjISNbTz9VVG4MpfEYkW8YzP+gAPvQdZPJom35yP8/pOIYgQIf+xnggvr1irdqEUZ0+ONhpUqqE
8b3L+OylzUYYeW1CiWSegOcaUNwEpohB1K4wyqF64UTfMtufcszKP/0VjhmLPPAhb6MLrEu3Y/Ud
0UmBg0bIVShxfLl/vM5apHkHkRUsWZ8OTExUq4Tu8bzGWgVMco6HUfEkCGamIA/N7uO+TcbQimcM
z5DwWF7dQUq4VaUFdAnrUZalmJxgyml6IwrZ5SwWlJaDOSUkFxXaZpVJYV9XX10q0yfCS4f1mKy+
MD0ZlpSkcQN215MGDE7bhi0yKwVNyRow4O1tn1XYLDUqCGgpncb5TaR7x4i/CA+LgDi7LpNMIw2c
cj0QTTUk0+PNFYxSAhrTBAEzidd/Oc1wgiZprqCmCLFIxM4jKthY+n/l4CbW0Hi1F9/vDh6oay8R
mmAUPAE/SX5615jg6P7kSYj2gQvYY84fUgJvBG6rGpm3YZYM8UAE+4txE5IfSbBswssgS3vSHddf
Set5hwqKqI8yHgRpR8Mu8h6vkO/NaLCIxAWaqNT0dSAGTVGoM9pfPKdDaSQVeTlSadwOFOOtthZn
y4U0ONUVNPKY88zWrVePZuFk6U8LdD8s6YQ7f8Hd0I2kWGOjEOyy4wmb0X3V7/OM+L3kG8Bl/XgA
atG+IQbxmxNEm5xnQDz3GCWIRE/v3P0G12PprACbz1UfLCENyevf3E/QN7ZfQxxeEtnxsDiJh/yg
6i0wMf+e4VOZNaEZMQJhzRyb2xSaiZnumNWCTxhIWfSSZ+t1FQFc0GQO58AAPxsUKYfEf8U77HIA
Twh1odKwU0EN7sFBA5kNLHISaHqG5KpgWvEqq9STeFAsSh4ZCLnuhnm8NVnA7zOkwynFCRda6Zzr
Tfxkn3VhLaDgZb34gYQgy/b2Z0MNNZ9Wa4dhFAzDdqKUBmHdtgBOQkVMX41/jJf+5TyGmqGgeIc5
OMsX5h+nYwkTImoBdmzvIAj/BbrbMq6mMomt2GvAFk+fDQUt3WcF+DLsuLsxZQL4Q5eai8xW/pmK
Fi/Z9ei5X18kX6rvpPHbTPX/+4A6hvX3kZgUulbKx5jSGOMpoccO79K+yRHRbczvBFEknmDAAZQM
1ZubdC4glfdG219YNkJV1C1K75lj7VsVd83Q7FFVbZ6Xr/DCBd1Npgey5b3UjrJnP22gsccwpw5L
GjV1FRQeyRb53LXpDjdefimQBfoCdQnChextolBZl8az7DEK0vgBSx2pDbHFSx90XO4umFwEZSQz
jydgQRY1tuJFIk01F2FteWVwCsYv2Q/3kVeu3tXq9QA+D39C+++MfoQUNxmNWTL1ndxosfHyZz5n
5/shpLpA58YzM0+JsmvAy51dquYEFyYphgHW8k39m3cgLc9FMYbWW2nO6aQ/yxFWy7NRjvR/jMwm
EjzVb6Y55P+D3oA6yEP554n6FvLYhPN16IFxp/WTcS2VWqYZ517doJxlSSASB2rcR0kJLbcvAGiN
R4rNU6XcuFyhuPQtoyk2u7/u8S0Ms5H919hZGzIU3bnGwpY7O8nxOw6xeqJJRWGhzOXplMNPHHhV
3FFAaJmwu12UyfYTUNqAH63tQmNQk+UmRsrRoGIZIy0BomVgW2gSQqFoTcSl18ypBzJWIvfXHCjp
ImbUWPKwPLKAxcR0R2XyQHgHLpSyDI+BfQWloDVBZmgP0gv6Cd5pZFycUf17KI0hYnN+MMKc+nbc
Pb/+HZ7oUQuSG+fQNz4yeVG45rtPHn3690rtElgjg61velcEw0FCoTySkmMFrXStdSJBKlyK25/k
6b1d9tzdcQAOtdCMegw1IYeHEHzAGMMSl/OLM7CcheYWR5SJX9BRUZnmKdX7ifozYwRACPb4RNLM
U45KKVKHuflPeI6ZrQqBU8TeYSMr7iGrZiy1WNyLn1sjKa0ozbnS9gFiTsfLfkTiqCxPJ0L76jmV
r3xF2u25XIx6Sr/9EWD9fn3rCOgcZ99qjsqIwi8URRAOLR/E0BF3JBVzWw+AG5h3cUWexoO3ZrYk
ChvjQFZV0jHm8K2IhPoJ+1OHQz/vHCkGU27Xm7dR/NMadku0BGwVZBWlszhX7ojFbWWVfIzIf85H
ppzy7tYpHzPTxutpDcBkiu/FE77ydT5XkgOK14n640IEcDKYBIbwgkONTWlI7sWud/AJeSTvfKlP
088T9jfVbjksX02WMQmjusOewg9ZGiL5Lv6FGMW0d6j2Jxn7Qb1Ns5BBWJP+MZRVj4pYvIF3iqe+
Pm9WzCA+iygoG87gOKL93b5wTla4jgSZIiUbLeplCf76tlmA59/v8eGxBjDp2moozMEWs5Wlb/iC
LJde5nf5R6muGeBW4y4CyyRkRt9Zeou9UJMYgflSc6tAGsKAYdVyYt/yJzJM7/A3qQa+ibkeEz4V
d5jFZ3NYlm0Bd2A5eLJHDayjhEBlzXoorSt465NNeXvn0Ruxv8s7VonfCFDAqItq2CTgm6Z+rkCW
J5CIwHvNZtXyx2TBgIOiNd4itsG4rUtdWTDePFfdWa+qhBHSqZskivWeMR5BnnDMpxofTh5mjo76
l6T3k9NHng+/B8tIceC40coyrqH5GM5VXsOsE2n3PoT2O3cVSFwGZp7fBjC80j/9yaZ4Xy65VeBq
/J4vZaHRJypZYRDgJ5vOVHtMYH2s9Ft5WyymYL9bJ9aXa/ESjQtnJHkooJtoxGWfcmEb/Tz/cYeu
z+83tjXiswxrcAH0JRR13Um5YycFIF43HUVViJdhQPCBbViCCcxPDIBx9dlcBz/lWo/OXWTgZGEI
B3O7JkLsGZHuJpfgPArzlyljc5cN5W1b2vlFv7jm4c0Pfd2UzZygt5Jaq1xkFCJ+RwesOvrhVXC0
agxIcb1bt0TB6waSiCBI23iLjYEsJ59fLrD6O21KwDNTGVbCZg9vGg4nk3wzV7O3s+//OwCpXOO0
fvCtniaf1+cu3csBFizgZPDy7O1+OTVOvUhWsu8Um4iAcg8TcHGbkfUJSAlrrhxVm+G+PTkGdvIU
jkJYMhHQcOlLoHaI19Q8O9N9yKGGlj3HQL1GBHXelPtxtFZ0CqyZXZIP+mEM+/wpjfz2mCSj400l
wAtG8xk7FBXcKuwC+kMde8tpdIksHy6PoYAd7HO84VzEKtiSSXYu6RaOF9fPFzhHJk8fePla1G8K
3jmwG2BLh0jfkkbx0WMrdPYELq4m6If10MoOxWk6Z2yE61+Ki5CX7YVSWd/JLQ1zIXml+fWqeYhA
tCUhAXFAuNWRBv3JULLyXPr0nXjYUHb0I38PTzUaRhw15NBWjyZBhdZVFV3XZ7mCx0sjnQwMhq9O
ijyemiSZqUAzUQEcsCO9c4ymBODekiSOPSaesqhVwtMoGKElnxvcicHjaJTXSh+KpbLnLpO5IXg6
CruPxmY6fJQDe09aVlRkdTB9MsJBNeYQnOM5exmM4REDynRZo7ZQvBvjKzcc1sD2CaB8R8p1AARH
u0+t8cEdB+53nPrJiT3DHFl4E8qUaGCf9tkL26MP0bHj7H3X+YLHVkfLUxiQlTWgRoLoQrQI2NaA
JhFzn5bhodjEygyVqdaa/mUI6Sx3bXZtuup6x+oEcPNliTLVHWiwIHDsOmDRlXjcCAhXf975GvxF
gSxuUQ3IRDQ6raY1TPgBSustkSakDZX8IjjtQy2GEy4RFiASg7+dxiUFKFPymZm/3sDEC6WHLCfJ
nqw6s+7tFUSYemTaAkekjko2i2ksM0bcXJfd2DtjuOuozjehnb0z0z9uwuR/dW5TaxRneDiW0VA2
MAX/VAxHUCMz7J+iXj8ZLPdw1J0U8Q79SRSJrat4uC3vjrRMHSug5I9W2VU83B6PwFDAvQJIoGZ+
U1jUWFC8jP7TeZO8Zx+1EoLpyne/MBnK9/iqSxdOnIFrIdk5KhPK9S5Fz2xXSHKmTxNMojvYh8C5
CRjJ37kBXjBwIjNOqwsHzD//qnUPqLeGKRfRDn5tKIlpAdAFAE7LmwCNbW+aUejSN9OG8mD+D4to
GoZMTR+aUIQuDegJkpErH8IdqWmaKUfERWX6HOCIXXyeIX170nqrPO7GLH5VhaA10JQu+fzkScJU
A9thRHucM38MMFOjINREkoV97Mfyhn9hF5BLt3H1/GBRC1f2QGkPTwojg67pEvX72XQERliAYMJ2
1wmotx/UZhhhDt+OOPbj/zaDWB71Xb6gK2j9zmQZWHl6qGmxuO0Uox6dmcBmeLum2ox+FoFS/LH0
TAYg7jbPH+5uV/sntLy+ZaV3OjKdSIm0EKxuWwczD2A2UQU4m5sAuRhGuyClLuzqZChOSBeZm3Yw
ySJvHDpBksxpEnL0kSI4n/aUZa0VfspQY3AN8RLednAYJjNGZ83jAgafATnmO5tUbYyg3x2Z2N6U
X1llyd/SA4dk0WKbeN6TLxVZ3vT2HFmoAxmLcJRi1il4psbxxADpPUQGN4Uj4lCiT9dsqFgYvIIC
h85eofDwaWfKUzA32C1im/3qLsovZZDL18A4zCYtoK4afggCYbf1cJ2BL7zquyBYrGLyB84v8Pi6
23q12O2c6ZEjUFRAmKiTRqnZCHALcR+ZLduTOxJYiJaIVs8cfbo46h727u/FFzFM9FV0JMc5rwjr
efDaug0qq1C5sp5dgpENFbiqFCRBChxrX544xM4BYLKA+masn5rzdcJBKFHTu4iXnKzQ/dhaGjE/
mx/3EHzEZLNVrYUzjjxoPa0H7+q8wnDCujfNXu7QPNVignmaqrfARo3tF9+muf1DtGQpdQBISfnj
cM+xC2A8KO9CPqfWaubY1X3s73/Grnn+9py0rT0pws5PDRAImZVKJOH25W6RnGFji1f1VYHUqaft
Ip5ZGb3GFd5GP6Adb0lUXk+XFFk78eytUJ5Yq+NhmYsovKuxVDHwkj4VR16Ff1cVjKzYVZg8SVvg
/H7YBm+zk6pZpRsrqaX8YNF2V5lrjlMXQALT72uA8w0+s62gWydtj0PI7AXcmwcgmuWUE7VNX9UE
kh32a7JBoUYRNAMOCsIjd0ZsCbbWIY3XqBWuJ20tKaJY86+Y1zdSBh04LB136+iENdJclgXB+g+s
dfPfdHw1sM/tlEDEx/oj81/Er/37eOH6mb/j9e+VHqHRuwyJ2mP6JUp9Yd7lX9RNLNJcGXY+iXC6
JZVaRRgioeWYe4vCzbS9dqqm/bYG9BrR2v69B2Zqfv6rgjV0Y3Ib64KElmwZKhaYYIfIw1DUU/En
6bi2bb18QjStgRvlyTu2NDwtkmO7k/l3u8xSNI0NAeMz58PuzLLXRcDu0MaEdae2YmwTMBV4bLrD
jDlVyhKiDzZhPFV6WoPKIaaCgwzjY8efEpy25aT5Ev/PpAVxt9rYm4PcBOhh+Eb4OpPmhg5mJDgP
I1h0O6wuplrSHrdcMLOh4JnPvcihBbrLC4V7s3TZ5yVbTPEsXh0F6e4pECwpf9kLiZMMwsFBkddu
sPOyUIgl3yB0xbQCMAiOJG/IwEyEBrLy8XWK1GxB60d+7J44BX+hFxy/9X9S5Xz1eBcfuWW+n96m
X2LqE5NCp9kCturJIVvXjOV5ekcaoReL62S7GtGN5m41WNkVVHl5q7hax68qEEU0k+zgy9zHFYtq
fS5OxJ7kYPVPQeOKnMTvc5eaXsD5H2m6aYHnMw3lukQWRyDu59UlFhWDvML0DxxgSZYZpFauRmGU
3P7N2fwE+/4f+cowKGeAzmASXzOIPK4o8kWHTbIUVwQkhZLVHemwnIlA1oA9tDisZDSe/jWmBD/2
rcJnq30yGN+k7b5g5JVI/bTPZpuzfNgmxXQK/NaHpmeMT45Rwem0gFOvtVMv7eADvriW/qE3hMQF
k68Dexjy1vL+eiu1vz1ryV8K3C6H5+Yu/9s4ZQa7wr40qwDQLo3gijRsSCHOXhOE1mkeMQu8ceGA
FNRrDudkZiA3cc/EPKm9938U3ZbE3lNxqnaNbBNrbs5jQUn6lKAPeRF0u8FW+U1hpmJYhR1Mgobz
fUcbdNVgcpKGO/NJSmPhLiQbX9C6yj3NcQlX1Jjwhr/Z4pjerc3A0buMUOUQuEEF9VEcgrd3/Sn2
WqWW7OOgL5tmfzNjmXezE7bMwP4UPhmOfcTmN6A0msG6ssEtRlla9TKY1JWFb4pUFSxPNrHwCf7z
UqyHXGKK+jx2i1LlI3X44NIdD0GziZskAHQiSqjiqB+xEvHCWMzTiByzNB/UlLFhGgxlSsGTR+Qn
Wl/MzBKGgXayk89IUrc0MOpur4/zWG7VZMVcTe9oMGzrKEN3XsxiX7N/2Y5+Hgtx/3x5R+xj9N9W
J3dXLsqVQIjrHG31r/Xf113hKATVcqiywLXDUOloeJzyfgIQE+dIARPaaFtcPlTw7VwyLkGO5gJe
spm1ByKJJAX0nALx0SlfJXVUmZ/jdyN38C8+PXn/TFje27XUwKS0JWtw0HSHKFbIyMW6B7hGyWZ1
FDZ9YIEnhqrT5oepAQ2wg0cf+3WdI0zKZIytjXZN6bquemQuIi0WL8N+Z0qwOhKG2DIu+Y7gNsGl
WzaUvq2GalUI8wuquok+o8H0NTvVwG+LYnU/lvegwwPjm3DpZgt7b5DCejLM+JUS1+El1HX+eHNj
cO9YSSsjFd+/S77P4FqkhyoHX+ynDxUcLy/2SW8mJMMKUm0p+xSUivVNzFyjlS5nElXzvVRB7P16
HLNlsA66vaEiu6ePyeYK7Qg/D9x5zB88vA1JgkpCV8S38svHjvWQsaWd2vxjQtLBDvJGcgu8zxBq
cjIsmAWo2RqbvjSm/TuSjgMOuvYbIk60t3aZew9H391wtWVcMgrLUrNYqLhj+q6nfvIGEyDEIwQ2
y1lJVvUrE4UMNEKVakA/mSbYd9pwkEQvtaqYn5aIh3XdTxf1L2EWz1C4GTKOsvaDsm6KqBhkPGSz
82bipHaFNc/fxQ2DrDpPyD8Z032V52B/mexnOr+lBstcECiaFEGqKA96b+045T56ARhfoP3B7m2d
8si7vLk9gQDD1OkcFuZbg4WsQlnamTPgdnXdobuz8iF1htC4/9or7UW6aJq2XbqR0AAg3HW2nTj4
5BNhD7moty5Q2/FGGMVeLKadobNnVdC/zfonUN/tm8iKekfZgiS/ZAsHYkhT6rEq3vt6vwftpbBt
Lx5/FWsZ/zuiWwIspEEonn1GGeoyn5rL6rFNlHt3pNON80MFKyfkwVipBhfnqET78qg24xOMb0qz
ElOL51TfULyjwyWXX7jNHM1pUnwdEI4Nnb8mbjLD/2qJh/UKupXcv8/GtC+zlNwo++PAvxttIbB3
NuuhAl34kUJLruZ128hPcg+veRIQ+gyetMvcyoWYCAZfyEXBfjhdONDfoVO45c1TcOvfHEoh7mg+
XwqoNGylaocXXmJkkOFifj1d2sOyqigSp7ginfxpP1WW2SJP3S6cHHfDI7CLfQtDa/tJGoACVvXI
DhkAe8FYxX8makriaRkMkAGVXcJUDbLGnd6ZCB2GozaeXvF4c850QT6ONbZNL8nFApjcHyujuLzN
969w8ehXzTK+UzJ5zXYNPUcCExMJRkcbULmvIB869LfqPpP7IcOx6l6/nCV4fnLuuvc1g2IalugH
ox+j2y2OJPWLpcxsDgv33Fyj5/HQQW8QYP22CSThU/i1C4SIiWEQtS0tL517zgW1gmGWt9yKTFT9
92YcJu2mEXA6vY3OhKxY8PpcFWJ1wMdUYuTCNOqlZBy6/Wvq7YY2uZf2JrZDi5TzMpmIGDTe5nX7
nFa0hBlGz512NgAS7Fzelz+JECybmzIEJaHm9wDJcJukR2/Y79bxMrup11DKS5U+72bFZzMjeDKV
OfPCtjGA7BSBnjzLZhKN95i6OFzKMEf2OyTrHHo4PXwvJ7ngOntyeZlS2EjJoyG5WvgdIIx/L/34
X9gW5sLPtsr6sV7+bGtXPFnpMxGuHdy6hdAOyeyqVDfxE2SxZbtnsNtjTHnu69EETxam0xAFVdth
G3dfow4JKl6oyWxg5gis1dsM3j+3TA41DRFE4m5eQ3VIP9aJn6ipOQzTuKtHoVSFN8uCfPYY3Qxs
Q5rlkJkl5P/kGHXy+2Lw3X/MGdQE6Sx2aaf6yuF8kKxIZGgpsdMUyH9B2R7fXQW6Jk9u3SmQeqy7
mP8km1cLozCYGZEnZ6ZA4fzUSVAgvdjSfeJXAMMRbykfPc9YZ2bDb8c5y6RpAS3e/ynTgHcB7Q+k
Vi3WJ1JBLGkgGCWe+avaKW8h0D7r5OOXtMIpe0HmzmQsD8KfmjTxxrU1+ZjT+8iGCGPfeblBkCPz
/LxGJcXqRWHwD+ZgSImDarM64dAU1UawG/4x1PBqvuls94gX2eqE3ZEMy7F0/z7nJ0B+aisgdJYJ
odGqlgol3sRQlKzPDioFUjpO016HB5e1gWEGAH5hfGjTNDtCpRXUg6HV9sBY9P6Ls+oCf7TfByoD
eIO3GnHH5uVgxZTqwzyNXqTZoipAg9GU8Sd1H8ri+XqYCPzrz1U9oqx2GdxizM5EEEq/nEH8BnLO
+upOdNeREfwnEBRjm56IlOzxVWU0lbeKRctnPlPNrY4JgxEN6h31jKbWp4LyTSwbiLC2cl1MusOR
sh8egR9Sa9YVmVFeSlbqbzUld7mJIIspb7JTWFUab6ck0YGhALM8m4iT+xxKw6Of2DZouQXzrkxF
sKpF6TKimcdOAYWUGM1zvIRiRZBkAMLkrmmgrwQRBG+FIigP3KGe5iPbPudNoCSyO7ytFcG9QWRl
P8PW1aCo20HDIfyWPGaEy1tP8EAia/l3EEjQzGzHASaRYRyboI0mG3vz1NgamH2aDW3gW27oqkDN
Lz9NpJ2w39qymopHH8YU26Zb0PEzm7dT4baHaQrABoQWTTwwkqnaMdYGwk+FPtf8ENBpMUqYOZU/
j2J0tuYCtUiJq3mq2BPq/YI4+/oZcLGDxq5MbQq7qlt2qQ0U5WhMHzjJJ0GjhqhZE4crTrOz7WWu
k7GSoGgOuAMUyjnug5OnjnUOC+1dw3mgjYebFbisStr+9ePmycYVJR0K/+vmaQAnbBim4QBxjfEJ
X88OYdA14UjD9GPqWkcmhGaKuYofsq5t1DSneNS/WGVDEgBOD1Ltqg1ZHLjaSNBikvbg/3Zafymu
+usVe44t1iZNOJqEUd9smzYdOOZEZ/3vVIlxf7mdU41Y3Chwj3vyWmkoTGgnniX00CRiTj9ulzS8
HW/GUuwBwb6ujpAcHrgCbrwmU04dA/AYfL9zwZYXQHZzpsIfTBKeYUmqNoP98o3fzJGRhxOZo1qd
7AsswJ3Eby6eH5bIsiqoO5NElEnzXme1xyosYFdcSIj3TCJCpzYlDSsDb8gnbJTjzGTxRJBLF717
diTDJj+IEjUAMi6QKD9igCkEh3Ew7WnarmTEgzcJ9WrwdrdjngyBLAkZDPl23SVJpEQj5HK7w0vW
nw3DVUO94GwXSMukLffsUlgHnL3vMEQB0lvjncVssSUFmkLewkzvl1Sz/x3e+P9PAj/wv8xwvrRf
K9N2fclV0HDLx4ZMeILU79MmTKzPxcM+scxCl6DB/NgO/j35JOZyRMZ3sSYYlaYKpFPzF5kCTYl6
HX2f9F8qD2Fea8C0x2hwi7VG6LY58wowMJGDwW+q794/viE0OvqX5QyQmwle6q4MfuHMqQaVeq3h
ix6qAh8u46aY/XEteSpswSqB6OxZHxlXLf3MW/wb1jMCT47uo7X4IevT9orShhYb3UAyQbvUpU/c
WXr5wbTX+36rjI88FKWh00kTty6v6HPP/iXD7dnmeNpLN7YaFJrQEXI3IB7NFnJ9ZWhvbiN+5qEN
SVtQm9dWv75fm/z1yXFgp7PcB94/40+ismE74ROrSypgjUrJOVOWMMhrJ8sx1wrhvb5WRP53q3Yf
P/cwL8fTy/BDxxnLkV+389EOmUc8s+rw0I/PAuGIIkMGR5HTsn4/qrY6r0cZMrf9XTmKWnA5PNP1
mnLpSpQmKzXkV3A3VTLBvFZLaCn73llEh2Dvn0qGy7F+Yuaa8sBpalTOdOA7Y8CLh6GA1xu+OaNM
QyG+ryc/vazTVZo1vcFDIPV6lRKDRR0jci0r5tgmJXj9m+g4XmqHVMptHjExnp/2DVquY2MdhzVs
KNodESEShzV+NregsDzk82szimDuKghiZRiPwaGbr8fW/sdK/KcWuSoaQpurxDdkEEzsfalfEnI5
WOlZKvZqM1t3Xr3SrSueh3JCMT/MXRyts11BMlLzYDhlds4UiJ0b2CWTVAY1fWYF+WRzvicighGN
QrQabeZrO+LFODkP0uryWYJjTQerJaOrKLzfHyqJ3ioub/4BQCXjANuGWvD9P9PiHpIIag36xPwK
pkTIpj+bWS0Qvg0t1C2hSCEuLuduUkidMl9zbKt7D7Vv8Gc0O1lyttsTBrXTxq7FjQZivtu0PLE5
gXEpRgVCtFxvlSVlDalmNLGnGonWpvHZwFTpBNjqxssX4E/bcnnngtjbhmxW1dkVwY+X3rIrpzd/
N+6BggWTKxQBbFElBpR/IlNyj+WOiP8Qoh29xD6fZsYfMHIApRQFaxQSzGikkSpD8dliJpVKr1G+
tkaxMmJpaaC70EuR7YKN84XGp7Aoy4a4BEfN2nOCeMCPTbz1NQ17KXfhbAnnY/jmKa75nkLA0TiV
NLJRK1Z3GM1H7vRr1gjXJha/g0ORT666vcRwtLL0KblAzEzQSuIgH2Jtvljn+2zyhoLQMfP5lhur
LRtt8Xd0/dIkgpw78T1+YgV9fy4Zk8t1FJsFnveJCPeGPa64taV32W6HVMhjDsAWrTQJah/fX8Q2
v5F0pImH/4DMltXyJFij7JJmJovcI38Ynjg9i80JRK9FFscn1fS/VwJhTadjfuGtb0ijo3ZuT6bg
7v3XSG/9d/dc8o8b1MYOzgX+cuOkjD6pIhQ4znCzQeZKJtYOd6EcgGJKkmDHxFrlmlNdzrJzQ7my
l08Big1O3yfFnXefs3HIcDiuHNRhMuhTBCF2PJi7l0qeWGVZGGNAaUEQougLCEcyokPtmBMkoyCw
zBBDhzPosgI96fcCj2nuEMlj7WO6GocVWhEab8dEyFGF86IiQOVO7Us4N4bfrJ1YlIUPgeMavbMN
LCzxHAu01AX1NhHL24bmP1r3DIzAO22fdzoW1vu8wrtAQbDK0W4Q2OZ9/xHzqEM4CSQODnDpT2hI
iXBY+IgEIQvILQNzuyaGh5QPI5CUVdnvXH18jLt/mdU0Bcp/WTYCWBU+OtiRDrcktCplNkbrEN+T
aJNms2dW6x9uelbHELF0KW5V1SV9NlTPSTnZLoXJaKwxeL0zJ8dvxS+J+pgxxzFJxr7XHyFj0h0c
1q/1F3+nvIdlu3DioNyHlDm7eZMK/90W0B/j90PfvyfkIQig34nH5NDk4pzFLpjM/jfCAvE6MO4v
y8DYZ4ICRybrU343xHyK7ofmjTQzsW1c0Yh9dKJ4V3EtmHBnqDt+lPTsO3dv/0B41Biql9cgmM3y
GjuB3wh8ka4daaYd9jMqAKJEIoLE8l9GQIZTgNfEhB/3GZ+35K93fRl4sq3WplUqxoig4901sDMm
GEyqkS2av3fmtEzBAyZakKa6c+c9zudwndkW19FHzvYc++dUfDkM+DSTxGno91AAyGNH1rApcZv6
8j5O05c0tuZ1xYXWhIJlC9b7afGQhnxPLjeNkTYnmEkOdpMqdDWjLbWJy8XXbnQuc79VDs+Y2L+5
9vpRmxooRpzQnDI1vRrXH1IzGHiGbRPVMeGtCzM7YV5z9NnamiA0K+Q1X8lIlGTb75bnWZr0db7X
QqU9JiIG7EBmPLT1MKjP4P3rC9KSiKxMjQ2CEk8WPKaiwJG0QA4aRFjjnVnBY8iwxecSSGyo8xCN
pJi8rU6+j01UaO3TSy05i486w/iaXZzy134I7298UOcZRGvxjjpAyigyFhkzers1mHb2NVNr4hk6
OlzSLphhi8lnurVpveEAjrQOQ6trcc4iYIo4l0u71NcusKGClHMtMgznhlV7g3ZGmFdQ4bRpAQeu
9x/4+DDUUmg92NW5rDCLGw+annqkotFBNsEIbyvX3uPMrh+kgWx3J+OhY4U+bESttiS74Nctd+6K
mmG13n0G5KqqmNZ2adyacsea1UaywR0eNWOmI4JSbW/YN01RzvcN8T6CzYtG99Ot1Ne9qALlZFzI
g/zOVaKzK+TSZz+DJpXuOsKbv6abkWTpWfy9XOvfktBgxla6d0EuATl+cUMDQlOMtrLXVqj2heTo
s7pVRHBDYHsR3hCxARP92kjPXbzc5DwJRVIP/pt/xN9xPt5Q0mWblQ8Qsb1T7LlIkKK7t+PImvWP
hNNQ3gWasThZm5FFzuaCo8IhRq7Wb4upDfq0GB3x20P5OOhg79fvBKJSx1URIFSDVt4fYD5IDEyv
srhfRkoEsse5nv2CBJaDmNz6+kCtrqeyW+sKILyivUFV8t7fUFSnEMVBqekDROx4W1XwB4cQjsdC
P2sCfyWELXshW2DWtbSSj5/oSzxWIka9Klu0jnpDdjvu//itAyFstToN3pRZHpn/nrV1fnd9kwKQ
3j6hJtV+wQYaRKk+jGsuF+bTxqdXnO20NxNUZpqCzu7/DtTTGtBANDImQ8SOlJ44PM6F+odJUXM9
HMbLmHliERICQAN/7Puk/86U5JCXuq1+wUGgGT/Cr1Fj8Q4rmueAEO/q10XrzlprFBpOLvcppRif
dx8efj/0h8NfTqI6Emv/KG8kcDjKffAt3acTq3zETQlt4xKN29Pqx6XTze+sjpM6Tb6CUNW3Od3L
TXcKMc2USbD1ZvDomfhmDBGMa9dGhcsaNCE2rkbemwhpk8mH4iwzP+3xHTOgIOpdF6D3JpwVdPDO
FDEEzzqaehA9wmK1oJEo8Rz5/A8T6MRyh+LxlQo68qa6H7BtT95mikHqo9+GrRDwQDYJUqwbGoEr
LzDzm4kFSZoIU97esiwpAdF02+IDYlpALkTNFyTfQONZZapxpBGQoPmULsOJHTsVFpU4vUgJ4Knv
ALevhoc+b3O3nJFSwML4afqzDCEQp5VIyLxKqn039Wa6sm2sOHaK4qMIyh+Nan1cazz0i0TwHfOF
zZoXTMst13+XsCtmwtbPGgM5HrfN6o14NYJMA1KCATJOXZSOaSJXZH9wYdARn3d+Khu8WoJ8GFqT
8+fjZaQqRPyJym8vOYbk0MRim1mX8ZoObwlg9xmIGb6ujA/d9f+9wCyw+fipwrsRc87wOsE7tBvy
KgJqzf94Y8eAKdQxeLg/M6iZeUGjtkT9TcEr6mXuTLutZCm9ADqGhPccn8o4BQ8INNnRCpZSDShO
1OWD41PBlaW+F1mqigaNMYuHBAcCSopVdZT2X58qpxqzJBF4mTbOEP4k+F5//WKMUXZYcRY0kVjq
PlYr+QY2EVsNuQR+fa7GIPTVkgKh9O2A2L3xZFMDFSEX1b4H7ZMPBFwLMe55YhAdj9XXerCeCedp
MFpae5qaDfru5Z2wALY/bBHCpFAXp4V3uLvyGM9CIqqbvgNuAfKeJ8pnRfeJAU17MxA7nKEZz4xd
E966GfKxWFSXob9LHWn4KwFqh8nOkFnWiGj/lqFUwR2NM5xZXYYWeL2XqYn9dpJ1MbN2q9kE+7eb
VplwCPsb5oVYuAmzZfKn5LZTl6Jtt/kTy2ThEqz8lec6n1/3SMj82H08Sc8DD8NI/oKnzLx5wU/s
BK9DckmKDkeuMAg3E3WWe+c01HF2q210NjV/43BELeYDYFFwndKQjAWdWMY9veRuSTTWRq2rR6Nw
2glJqLD8JzPgwUOXsXQcPktd51beUSXSZm9cb51esyLsZqZ8bRadmnkLwSXGDJEGztfZfadso1sl
t/aMksTUVAPnUtfSUbZiDxHydSJ2+Up+SYL1dZieK7aGO3FqIT9yeReOxN+1CrrYUumdY2aSepx0
n2Kiqe+Ug/p8SFmX4mDlvSydJ6YVjNhUF3bO13WVzTwvX+YIOzfal/JevsdHEgrts6aBcqmYg1aW
EUQm3tHa0LQyoQXq4tlJcVIED4bLFi0NAbHg3/OhMiLzuhimqUOO4oWmKnMyF42BPvAbGi5e6myZ
bxv5z0p/Yu5Sxj1khJ6wGo9D7uCXPmD4HkMXXfH69nqbdkX2DZ016pCGVqEzfkOwD+BSqdYeNhvL
XbK9vIJIddjdOfqRKxP0Pz5HwJj2Dfg9MrBlHrli7mvNnsj4XgXRRKf+AJYBVw5vkdLj3mmGBh5K
ue6bUDIcQZCT47OttE+mpmQATwk2BMr85uBr9eyRQaUSbiNXuFwJ9v+DnW42e3O8LPqo705pIUSW
rSwxPjnuHR1ba8ED+DByYODu+Ivl4fnx9yDe4XDXf1VJLzQGojfUOkWS6o8/0qd6p9agF2M0LQnS
mzgEno3zHYuz+4kBAqiHDsZ1ppOzhWX40wNf3327SFLm6H9bbTaex2gFUWUhHm/OrN1PXbaiCcQa
FdlPZYJ51Joro5b4OQEWDet7vk1rOweatZcYGpELgGazNfC5r7ms7IQktSZiSfQVWVnZsm0gJvdi
DvgiXSJGGPA4qVF/EoIP2z/NQ3Q8JPw2P7laoqybLhM0m9IWRqPZcoCdQp+7rXhdwq6yVVnei35W
xwEC31t2oJiyaB0nosN8BALCw28LSIUv/eS7hqDOJ2sB8J+Y6yeCn+oJ31uwxEuN2KYCfqdhpoiZ
EfLK5aUWDku2NMKyVHPBkr28hkbFHEks0R3tq+9ubriGYd/FRzz/+acnwfArf+8T/akHD09p8hm1
Ox6DMF5We3xcgDqkVvUa2Sq1l2tVmNYSWpux3BpkHc/0zv+Ufl3jJgAQrBIKWqg5ifOEelQ8scs5
5U6bsm8OrEdkYWPDNtuwjMEsn8VVdsgy+YWc2Y1tdziyt7LLB4ImTuVdwv7xW/5Gi+gas+2rPMjR
maS5cmRX+CYVAyQZm79a/1nRUr8xpaGQQq59At4LcKVWRKdlgcY0KGUyYHzN4ixvjkEDE6MbflIg
fw6DPo0ZlYRAFTfXj6AfZGvTPlfScD5RZrknRtrSjyRnAYtbvPvdebv0BfihAFhafaKZVMQxMOd1
FIw3nuXpkyfVdwlMiDH2zbwE7PuE16jqMs1/3WZzOcP4rB+Kvjej5wBf70Cs+dmJZRpOreJ6wbHZ
kphx5/9WkRzQEgzImFVDjAT+FzsyqsN9hC3AdBd4ImNqr2E/1Up8khFeQOFHLVcITzNQK8okTzBo
vkhGVMugRBVCOjhRwE37lvQtNmUNJ+6plQkLkgH87G46dFQklMYVSTasSEPCcCG3IBHlEa1dNtgV
QkYFD2+BEddIFV7Rfiw/840Dhm+CrzTTC2dhduBZ4g64TgEXdSyX1MM/QPL50LxtaQnS+s1ylvie
cr8mpmR/IFkHmbtzwpcyUKswHGn0gvjDqmNwcA/hjNnXARyhXiFF1S5aV+WYuBHjNYQPlgzUCI/S
D4cljk5IsZph3WJxy0acjvD8qWKbw6Nnyp+ZRdRcxm4nM8F+QdjoQHznkHL+GJR5R4Q3QXyP2BJ5
J4X2/5IZAnnDesI8LZs5xNv1GM4HbbOQhnkwCqYCn0A64imb2X++1hwcVDk1h9GWONVqodepNkE+
qK4150Ag9R1ngyL02g/bkOD8/LsVXJFDa5wgp13eN47Imk3LGfl7/t2SvwogBd3aBpFPXYSnue36
mq64vVk1bSrMM3bt9JyjUFXpvTIqXFT/RHqZ3teRfgmcz9JnhBsZqQVdKP0ivaDtiHBGx09HNB2R
85wAyPqjx0/CygTfwIiX72e4NC9hB0kRsFHy7rzU4wxcMsCxgTsOL/2UTx5Qu29JuNJ+pqvKvLTW
upaU+3BvUSqnokbZtOWopq+773/5Ud/jsd6vKCyW1YxCCDCwYHDHbtcX5ZDf0JFp/bZRXT2Gs+MJ
eSFWR0gYCSPRsE3MA2e5wtlN/TewtxB1htFagrMBsHXTMiiqRjgSL5/X+TrIpMp5nwpmbSTtxQb5
eN+phTaxD/EjdWvt1ZZLpyMV8Q3W7KnAm7asfi+IUvjX/Qb3OpNLYzQKlXerTu0Y81w8kws+RHQq
WzKSNEAKL0kUyGr9Ovk8xGJJrdWGT/+8SYJZVhn2iTJU/c7m0i/XiqA4XvGQMWmSddVxPA7hsmFa
081I4Cu/XU8If6ZSeZ/DkwkYer9gwvnShHgrOf0+MqMdSX9txGQOtnhVUVaS4oZrgAvbn7MhxBgH
BLswRT80mljGS/1oKEc81XYLkGItXIeBAAsQToHwjK+VdYb/vItBmXnKCl6cibsSzr0LS9ANGCL8
a0DA2TF5C0YsmTQO6hcgUAsBrrDhv2lqB9A2H6joONxZL05UWkZlY+QA961AStK0x1SkjCAOvMcp
oRiySYp2JYrj9hy6tEUGJBGhH9LiP71GzSolAntNVHyNyizZ+JNWDTyaZ8zuuBW2BZFF7YUCC5ZM
pzrQUljLs7G5duFzOxJT2YyBzRn3o1Yrg7gMvUV4jpLEXy30hJ90SxwOsP3GyElilLn2UxbVkCdU
Dqc91ZV9Zbnr1JrpSRsz6WPvU+RNey6HpDiNUaZ6OfcG3IN78bs6pbllZmdUQtbry4o6gUfN/FP1
eAekmHMj5z/LMUmCLbtM+hKKdjjZSLZqFgD9kb0ymO+rn3xKDfX1UEREo1ucj/X1QzJvTAnqVEQC
sdPvW/bpJwPLcPyWw2QIMcinypvgTiXZ7qaHF53VV6UgWYKbSdCvNuV/mTF0lbvCw9EHyFsLBH15
cjTkx/uoVCQbl7pty8SdvGkuA9P3bpbp5jCuqLMTFIyIU/Pl082+5nR0CQNvQ3FvgRZMBCwWTRAH
sZvBmtShV2iyxU2JVegMokKTT0qFGPwk9YEgqlFFVF6WS5nOj//8W4sIbLJ0hajVyEPZxrNwE5F5
Q4ovVjhC65Loa9c7GYk6YA070+FqZ8/Xmu0IRlZhCnWs7DyJCFdPKuBbxEBng7eXbyBqdrOWGoBL
W5U8PgYxPAAK1P8Rz44QcGEFP43Ac7FCXPE8Cdv8rDecVsvAdRldnjqFrHfkZeZmaqIeMuzFOBBq
p7I/X3+icpolJP1/VKeG8ek6+8vmwm/gW/KpTS18Oc0CghGyM40rww6F+jTt2Zw864TjxMoLC79L
FNLUFaus6ByZBWYrBecMi7ZHBxg8+ehBF4KPDcZ0B3Fg5fa8b92kwEjYqMCnHT4u8Y97pqvwYT7B
nfJ7ZL3F4xJFjKJv+Bk4nQLQtXaaNN0JSgR80jCisf419kNb2G8L04M52DnVPglgigbiTs9ceSkY
qBuGEwWScgzCDP1AzwrXlIQFrRbe/wfgTgceKMdGgE8CuCB6cvRa1HjCgHhgWkryjTbFERYTNXiv
ScRECbkRUJr9/liX4ga/WszzD1Mogroxie5E9dcXzL9u624U9UbF1+eJ36daicKj2NyrIkppwOJb
MoZ7aD1bkkVqxNLIfc+kYlvlCoAOPbC2JaWmIjrCvoGa42l1oyjjOBwAy9M/TyYPH6tdSgx6/LcB
+KPABj5eGcrx+c0t5yk2T1gqPDf5YQnUwxdcgKweq6RtRt+vHoC2C7iR80YYPXBfcmJUYepoGmJm
yUNt2k6CORpI/uIGjmLT0CpMZ20SWsJlEwch9D34mX2BrIiaGdiMn8jnqvWU3UbWwXafA1HTfm60
6Z4ytqgYOVQkEtp9UQMK6mYqvkqz6pkSlh1xHQg2Vrpti8ELZfiOam5UbEqR/Q3EjlfeVNbXLep7
EynWVEW8SehhSKPkBev4q3+ecjWs6f5tIPTmfqqOiFt5eJqL+8USwDPGTuZsSBOuJxYqsiC4LlVO
p1NqprQUHTCmSkpyv20UfXdnzHrjw3xn5QsGAMNV880chz27ykOJnTROICvu83Gu3Ap1FM+jBYDC
A7UNlmHgyqkMDFStuynlK/Og9uXnE1WrJPu9GAsDgDFNonbXY4cDOkWEyEGf/nsfwodiZbDMEjTN
h6wa+qM2xFHW7qP8Nqzi3lEYOGXrnA1qgstr1d31cSiNoxE19nbZ5ENJy7uXT2vujPFAlOmIz/iB
/5hw0btyA2GdyBhVq1GeovlGlZOqJqcU56+/XP2h7TGU51cQWFDb9kZIAR3/iRmjku930VLvgupG
Zezcg+p19IA8Qqq7LGyNZJND8UwOEeq1H6pUlX+XIWzgNC0adICriJkvZ/8uwTQA9fH3RZuQ7Awy
qa7Qebd1w+qeqWaLRB+kpGdpPPi4ud3B4MEyKm+VuwGLXohsCquIBU+SNS+6OWnZMkZN/hn8PHkr
Y3XB/99lme3O0H3xVOamS3mnP6Qrt1xFm072fHiJyqP5ZOn7RyazMovXX86eUygjcuPe7kijAR4m
C7IkBriCceatEH8zQc0pwKtn3S8F0JvT32tXVmyl1U3BiC1/pGQOizYwU3vZgPyzAlftJzEjWxpT
MUiLZuBORMmFRdjxWDDg67F4ZZ32qF661uJkT82gn4JWJ19/cnZxYCh4sW/O0HHFDjZhqkQfLnmv
wahnGcEgCc/FkQTE0HjepdFd1L3QMPjLBdF5QkM7hTAM4PAGkLqYInHAJVDCwqfssqz7zbMsi7px
yF61Z/vRCP+h5Sy+HLgIVNRIQAziq22BKU3lTZxgJ3rNcykJdnemlIdm7tE0FHNqm7quQXeS+b7T
7cosu00/j+ehZdmFiLQJuIzVj+4s/Kw8qgFa0IDGQdMsXAHPqMkyitkzE74lB6PN0kUSfM/crFLY
K9T5MvVfJhch4A0UYyy2nxN/EorWOun/IAwfCdvFv2/ySIvDMxS6aPeIe283Hjm34oo3yfg0KnDr
bk3tg2cVQwdWhTtasQgmDF5ctCulfJkF/Xo9yC8bVU+lBJuSF5sn5cRrNLeOxV27ZpJdo5dR54YD
UI+LWMcR5feBNLm437Rx1EQ4uDlWq9wUxM47tUafR+zRUqGL0ZXRr5054NDraVZ0Vm3WldG4dLnu
EddbAVuLPBJIVjQSWmJYYJoPXxZR8muE2iPCjvObRzv80MK0L8ld2hjp1w2ExQg+wlMGuGDYkrsq
8R3yFmIZo5ii6yuu4zS+5fPtqmOabv84S4g31hUgi2FTihWBtaFz2rSrLczGC4pE28wHtiGlWW2r
m7ZAu8nwR7KrWv9Qgw2u/muSoyVrZSuPrFNq91qoF3ktxSKYrKILSKAz59NHpZlM6qJGXOpCtZdd
D6wLaWikCZdJJjXJvaRUfcj1/sqmbAjbz+bK/5U+Qn+Frl3Rw/cXg5X6upv0Wjv/D3zN/4R7MDzJ
PyAO8zqPwnF2YoqC9CzzwlBZInwBSRu0SAO0Tox50FAnkmISeEornrFSF2bZMQxlUsz2oPp+1+7X
C8ciIYQAUS3muC5bBgSSFv42KP3SPfsHNAwDhNYPjYjeTi1MHU5Kc9R8+iL0EuVy4j+LDBZ1fa1U
QQEnO5gb7L7MjEGYljHqMwg9285s0psNDuqBppcmloTKyUOmDrCqCzqOHNXJUNEOGVZTvlzc+D39
4e4vqV79uKGi5r2lBFy+nGwVshRYfDtuLuuCRQ6+1LqVuF87w4Qjp9iWEHP3v7AURd+QZHLDwXBU
3B7Tc8ZfxwFFvUl0Gq2Hnpw8S21JHtnqGEX/DvJ2a8oTmreQUc1JhK1iEBioYdO5Y0f6ofj9w3ct
FqEbwmg+/M9hq7Ci3lft4Yoq6BuiUFDc5DaWs0ji79ttxJRjGbdukBLCA86JKp3saAD2UMItFRKi
Lboxe+mOGR+HDgl31ueIAoRaDGsFGCV5Tz7tX7K3AqiLBXurk/Xvpv24hH9uijpj5EGvQwZbsF2M
lLwaFnvi1HJE7rk6r/p2+x/ohrwhTOuoFElXMsNrbfB5AdHiw9JBZjeiLeatQIeh6etO591sLyQU
IiX288xRnCqr8dKiyMb1FXMUi1DHsa0OZF57qXmTBObzlh5MwqUQc1ugYldbrFqaqIBNy12Ze3FC
UOCcGwNk3CJmIO5dkf4EQvBKkov8Tn8k/D3O6DttVYYCzCgT7XD3+jvzqMVI6pDIhe72lDH3SZEX
ys1XHp3dABSD9HwrViUn9c2jh0UXu/A/rHYlXlJBORng/r1fuuJHMUU/xrCkgmyU/wFdX4Vg10fX
FH2AVlY9H98tSeIYP+V3ldzLkTVCeQJNeBuMjiOI6Gen47rcjQLMhxTtg8fVhZDj3h16TxzMwxhE
GZz6VNkHzIRwqSjZZEGw1n9glbQZdObAe6Y/d323KJPhmduAXX+gpv/KmxHXgzzsRD7E1hJ22B7o
SYnyjYQixQd4Nz9skXTXhW4xkWzhxqyXO46NZwa0FhadG28WSDpNRdc8//8qw34auIQqNj2iytb+
MoAj+OMOTC/NoZd3XQW6SaTVEi6Fkzp2yWp6HSlCYnXFXNuUcCG0aSR5Kdob4h1JmGFRfQdUHLSL
ZUqe/x66CSaaAEVQ3uuucKI8jWhhq/6r6tdpkccWfmoxEKH6wif3zDGr4U1hsoPlbnc5RLkm7mgw
j3fYJNNxPncUIzBfFVaR0COQbK8r1TAj0rE2e7MgxX0fmvOzX8fvjxxP8EDzVBworNiEAIxo/qij
Yue/kPx/9WA/vKFxjFegveWSvqeaZjPZ8xPdXLPBm5SHiH4SQYFWSnDW+r85NWnxq3vPFRQPhN5m
5epVBT7m2ACtlweeF/VBDyE/nn9RgHK/Y2GOKjuz9KUS7xWwa9a1WF/+WaATdRZV0wtg49W5qNFD
BxcphpP0Pw69ZCptfcHZqFWaJpkXLWHVj/otjMDlS2d4VkgBOxwvGhcDo907hN9uL2WGuKuE4/hJ
J6PKrqxA32y0BJpgh6lxiCPfRfXRUdyZXjDrpN6wFbpmQ2+B62+4pgP8Q2cZa4mRzRfMamsU6z0w
7r1ilP+lfJvpeFk3/9uQjCl8dSDvFgnU+fWgMMTeRozMvOuvq0FlXP+v6NWHukKIuOAfPk9F9C1w
L3uXbf5WxEdM5ye4UY0eOFUVwy8r3wR+LgR3drnE/cYG5H6R9CDQ/o9TqZkKSh1VyA8gy8WPrDhn
Inoal5kuHTlNXg13QlqAQnjBBncfb18vkynHfdgmaSk1K6Pi5cuFR1asUAMWuiSIU4wIZNRnRFpE
YeFMG5NbR3UKvqiu5uWuZsgmB1lC5C++04RQhpSIgvHQKthVPSadjZKeiMIJZ6tzZRSPsN3SyyST
g6yRr1wZixdX74bFKnAqwcuicZpZD+XmvcQwxkacnaQdq3T0ChZaXUdWYJomWdBOEbR1r/nnu4ff
24WJpikA6GySBJPCwBPeaB5mwMRRtASV723HkWsl0jzbWxdzKreg2EVlhfxU1//krl9E+gzUH+Wt
VS92T2bU2Q4krRneaiLhudKYzRpK1NZr9nd7J24GO0T2vJm7bGrjZcfUaSkbLzM0UAtpZyYrnqsj
D6JzvqX7L27l/VAlT9Wfr8Xl1uYGMzU/g7seXsmBFC4UHHUc079zvHCV1cR5Tjn3W92XxAOaBTqu
SA8WLftGsaCw3LtIfdiJkD0SE/ATJHZ+6WlUaftzGwvAc6zsD641B+RUK2Yuc0TubeJYPZjlLtVF
+ZSSFDn8kfx6mA2IvTmDJALh86zWJpi8s7rWwMeF4OPyAbv694uA7ITa3pfxr0W8jr3Gac0/6WN/
7PG4Mr6XdFlQIUyiLfYHLAGWUOnwfCyPDeMVaT8zkEsQmdY8CD/lQzOq10EX65FI7Rz6KyorFVlL
HIRWFCBuvuhSZ4iDRZg0ugH43PO9omiKfCS/iSsJksmITg8ppWZG9bQ8vX4TDA524cXr9+mUyqfT
jdlFu/PhKliXCQpUotBn/aZD7wbH/gM/GuebeMPLtpAAStjID7NXpVqasvPNExjMV1YyXotVfRYY
CdZJ6+G5+iyeIxgvf6M8fKnGrlpi3yTOOpxdytuq0jAQK0qgFEslVhn/LeC4gI40FcjhO/TQtKBE
e77H5BScfBwSGHH7aKwMVkmRacpOLtxm7ba+wzKL2ZcufIkrTmLMMYwkPHKnQCi2mFNLT8XjgpSB
jPJjH3gdZvXl7S6OyTjiyHOuSo8RmqXQ2DjvPCxEU/C7IhhgNKzn8MaaRKfhd9Fl+vV/oEp4aqeO
Z5r7vGrDsFTIKIRLIoLCavCs//T+L1N08kWV0twkWsP+K7G4zZFDvC42Tt0dYt7KHamqD3e/4M6i
f/MXh5s1XPo/XRNHXWtBTT1E5FH39kGfparS/q0RyaJ+3sWmnL+tId8EdFUwrmk7eN2Ipaqe4t36
dJTsWbkkwew7vvyY8jU0zGzAQPM1WADo7Srz0IwGSAOklSoW7R+oyMkTwBsDj7fxA3qagBN6hdRe
nGFT8qgNMUui6vdPeK273xTypEemA451VE6W2HY2iKMmK35vjhhWy0fkm2z2mlKzaihHQLORntqq
QKkWr+QoyvFy7OYPR1njR3BdfUd4F8nRtTKo8K5asXJ+O9axwRrJxf1uC+vbMqdioX5147z1P1rH
6J8Qub5iea32sH7uyRaio550eZs1EQI0S8A5ZpJQNYdDA1JUFWtubLK7eW95Ax7VOY9xEvSkplPp
L/pmGACf1A87zLxmL2O34ELckjqprICa0yjIlkpogWrG47LzeQQ102Q3Ai1NL0Xek5C8J/2s/h6H
k0tmYh0jCfi6JHBwXfZ8edP8UzYPbpDQo4lvEHtgyjhV6C+Z+uxWo5mPylk+/3aD6uyvp4rSf1Ea
FWbhGyMGkllOxckPzdSCJkz2RX4H6L4ic+gEln/iZ0JOUUs3VeyObUms4tDFHpYenrDJXSnTiqNk
DvAu3fKjh1/KQyxZKTgKbp0Rt2S+Ow5ddQ80KYEdGQ5ZW7u/ssnF2P3wfdxpeDthipMs++ZeyfOT
Mz8fNlIfGmEvma/odaKknUOmMw3xlfjr6bosNs82Qk+QWNgWzftoIuHNwX8shYWok59oensU7NPY
EN1YjYZrjlbv/QW/PuEsiaVKL99MjJKkdfcPyHZ1Qhq53Ia+UdnDBkaKFETBRbRt7kVDH6n/Awyj
4l2Ay8RU62MP97bky/Jmw//swC1pqQ3okw2AdA9ihjrvvMuFjfSSeN/IkDy04MEQ95/63gaF5JX7
mkA10vi6R1TRsaVQwXVn+Pp0tRpPf5V5UY6vhJ3DqHQmS/zs11hQS4gb+k6rvdWuIwrURkebtsmm
m1RUygcMjEVFVp3mDFVSbhI/2i/+IFB+bXyfx0zPoq0+DkFzhAS+94DCwdERTpUFbwmVXkSI9n/o
QwgrLQHzN4X0TkoXWJjcjy+X05AeHH1hMVEh4rrID5/7owlEJTJ85qRn1d8fYWVBNmrO/Wyk3btB
6/hEW78Um4mcJ+LPF2hGPX/+SSSRaSnW0NEdKZjCJSM8nHra+rByvmy1vYn737sQ0OM4bb0xTLAf
KS54tZnEL7kl5i70JOqv6hKS93mxc46r07CIyd06tngYwWYWWENRXmX2kUKaG5Rxd9cZTLFVHDWm
DAqtlcs7y2P+FImvq+5gqYLcfQnQu4bKwdToxHLG5DptA91lXhLg+nzJ6OR3xaperXaAbrRp1Bht
HuTn6uHu1Xpubv3pfEsk4MljFfKNIb5XruP02Njq2KDsmiFk7eaXuINOVH6wn46WH0WkW5Xs01d8
LglO92/ZfysU6ZyNYkMiS74TQSCzAox6p06h/gk61zwEibbQLLlB3JBAdX0+aP+NrGe0ywLCwB60
T41TcF9LZtSnbIU9P+qIq1wab+xL+r671EwbW0jgFNL8Q0lEwfMfjtRI9aPDJ5HE7jwm0wCAORxt
wBBKzKsQjgIqLlfUdSohNalp4IAbHxXohAVb0QmOSZcw8/ifpMzEPrRMm8EEevLN9c8es4XO1ErJ
K1o2E8TiAKRyAU/RbJvn99zB8KxqjVZm0IAEpq5meUHNTCIazi6qwZFaK/jSgA6BcVf2ngf8YMvj
04CyYS9N0fgJNDZuy+Y/Jnj7DJAUgcX0dRa50ZjcVLcN7QvsGGn2iM6IlSjhcusTBq4F9lGnsxKn
KdJMrjy1aJrRx3nRqIBKaeJOf4mDC4i8mis0ej6kHzEE/WCmrgjU1r8KSZqmx+4DmWZxUGs8gxOE
W1izdH5C86lyUHjDKq1U478ovj9Wm/tqwyEZkrEY6zuaeAWAvioVGRM5xXBSHn0n6Ba3EtUl1T28
r5Rk6V+Wu2gSkEIi5lKjBt7Q//QFDjtb9MpJsNY6CyzhSMaYB1wL96F3C+F8lpT/R6w+3lTz/DTu
sG1P28PRj4KbjirLUffYCUAufc33g2E0nrzLM9as1+7f+IO2gPPp07KRc1z7NleIlF1gEC+MHoj7
DNo//2LA6qp2h7eCobBPCoAukslcYf0F7VXwpXSUbYzwtgJp72GdVTYKFanDiflktWkqIo3SVNqN
5wBvDd6axBRk4FXx5zHbXEdZLbDjblNpotTjpLbA6D38fTt3rL/tSXv/M3doxUed2WJ8h2pJ0uDy
BrU5gfUg/E9xYK1sDwtnMBXMx0GRC69rbdzWCiJgiB5RpqlByD/IRPD+JL2PxB1W5pxu/jiMQWgM
N6trFC2gxSJh8bBIT6VnDHvQsETnvDl4Vu2TNO1+KOcp/arL8Uhrk13AoNNgUvDegXy/v1oVavYG
n3mqNPFwe7yWf8dKHEygLC65kLQlYLgr1snLki5uKYSjcxO8/8JLYy58/f5O59xwvHB87PyKhOpo
hiKyb4XwC3jtgXEoqE9Kbd0ysuaSazxhOCikCULW9l20KDk+mkqGOBxGndBV+tMsvKy4PMhZ+uUr
AgL3EQ5QEyNftt4ttpzI31zgfJRtgt0DCW3S+SCzIcdDdD6/VXh2Fhps/88SUv5FNLgupwiq138T
oqRqzXnL0VXHZXmQSIb2/hYEBgvMnmDr7rVTsuxgGh/ijD4OYwNzIHRjZ4vj5Mc95tPuttTESh2V
DqNpJYkEWBQMYFkfCyVO0YY4vgEtbdoCbQY2wFiC+SCrqGuQnvOiDUZzhMUgCiXYIpHzYUfA1QFK
2olETt4RM1Rv8DbViLCsCN//zP2Bd9gylVEQEZv3S8RIHs0dWw4wFdkfbgZJ/wsL9q3S8OtLZcUp
WGwVaRuvK4P1cCU6Q7jJr6+6zxFGoaveH9bRlUaNVRG9Pt9fU584vsQt/8G0IsqGGW7YNBZcjZsA
+HTDp0iJrsNtiOoFz9cLrPpzy9BtT7jl3VSRAzkgnH+Ln58sm0jTVift5I9f162ZmJfoc9tsq2EF
qLWGYWTA25iZtoI9NvfCl+aB2T2br7aQviRvnWFgzJSIzXUZ+Z/mo6BXsn/43Ts/0oFSwt1Za/49
bOPaBHZyV9SS7zBqd5cWC+4EgOJNbh4G1drSC3WGC7wrKOjYArL+0GJUbIq8ifcEhNHpyjvhsYdT
SJg/aB+Snuc/YJcALVfAN3k21PmUIAdkweWHhAIOvMsel7RCjZTuhojn9s8ROFj3P3e9tJnNQQZk
bu+0HO2WiXtOXRuT1jiAj0rSIBS2FOIAPOEGH/e3Szr2A4TqC655zd3YpG/NJd4xOTqRb153GIWs
XySj97Q2vsTyxNFDnQ24yRBd9VzJMjprzLyON+6PEb+XJbshyqZi8D87Eq3geVgvfok2sumEmrc2
DlyaxiVvo65VPWzZ0KEEld9HXszixpDH3c3RW+X+KhalfN0uFDOusmHJhkr7Fx8hBMriC5rteSSn
dnTefP9RIYsoL2/07BfEBSbZB2hXeY16CjQnX4gyUTCOXz9nhjU1mCY0ySua/80yNJcIPedp26/J
SYiUIhR75e48t7u5dOSKYTbRIJ7znilVK6wVevTIIFf+uXMUsmdL9UgfeRWQRoA3RxGRKEqeRNLD
T2niWSeY5kOLHzAZrPis/oRhABF17V+4+M2taVs/H1tS+5ZcCMFTal26DZjCEH7QlGMEepaLKGAT
sPhGjw+GNGoXZMFJlJSuXaZJgdhNEzpr0WDg/YXwxiHPsWH4dCMv5mCycYloKFWI/dkbxXqpxfDh
Ho30FPyFnev56/daHJ9l5jGZvkJHnhSEOYGJDVmbVIcixQ3IJXxfYrVYnQFCtiWcoNtvrWuEQKHW
R1dgQ35BdCjuXqe/KR/X62sUfalBDdohKIgD8GKQxCTU5Aai01cCORlv6MBKEebT2sgILW3m7wcS
JL6/LW0tW16N7BrQ62VTg5AdJgIYZG2c7vQcfoKnDHOVagIqj53e+JU7FAto+nVO/NiWinQOqYCw
lAhoPJV9gtCRb9rag9fAULMb89UEKOD7i0sk7cbIIAiNqChmVuDAQR76Jwx9lV1JsTgcWL959JXS
IG8/9Qalrf350L/i54XjbtWuNaOG1OkdPbuGTyzHuLEyckXeUNehG2zzP+6yowcseOMwJycksO52
EWbtGZ2325oSVhqFhsNNQ6Hr9QOL0r8POK6KAHElrRTPnshhl00l5PGwJQxYOelPbFM9RclrSov1
IuXnzXbt3VVu1ylm789qrHBaXUZhmJav4XUTF6nXDAR+vkYi7KAE4v6CWbJSM5LA8wTh7dy7th0t
qdHAvZi7mwdKPy3hmw+CfcGfdROUUbIupezYzGNXVWvErTVQtdMrZu4t9FrjhEOKXJKWzqbvKTdf
t/tlLM8FNI1CUN9TKCtAgsN82oW/+FED/HMZLkuWOg9009NqeombYKZ6IOf3B0gx7yyfgZlFDoH8
dEir2J8N5FruT+EKi0HeF9AnTI8kG2O4GRmQow95PFM+vjFuDdZOmuIxDBuWPGVO/dvCi0ohuILp
Jx4LiMiYsY2xG2O8HfN9BJ6CB44pkIZO/StEeXARDEj6NjQnmi2o3jRE2unqde9xyfh+sw/StMBf
c8bRfrWLNtdHIoTYhMLZM9X33rvBAvwxwKz4RMnFazI1e4DbUxMc/niQDHwgU8hvcqgZ4LeBISEJ
LMf4LvUTBcNurgecymI+KnBUlYsYEhcYyxqXE1jNoO+AlOyU+mo7eYpU828VqOVB99hTTwbSaeSt
Qqb4B4oOFR0s8pA8QkQcuP/dwL0oYCOCct6EUJ2FhMpwi2XokhdBQpHVgAdi0bv8qEgP+69QrAhp
W9y+H63/ZLjXGQXWTceBi4C9877+oZdvGORXwXL7bLnl+qA7IdZGv5svo05Af8OoTnTkBz/5DCpb
K2S5LY0yTiZvggtMNboAbbbJ7g3o59kCGGE1eN7jmHiySWMhkhu05HcrQg8nuTX5SNnGeridvU5S
T8ICzTSOeTvuG4djVgZ5b8dGSYvCd+NrvXB0QgcImjNf00stfelgy5enKpyf+uutB+Yc4ncsSZhk
fYVc44i01cJvBbXpcgSQZprEinFlc8NElQcL/PBe3uLdrZI5wxdCD1Rkoaz2l0RlNZLbSJ+21CYj
vZfINvO5slS3PgsSFRrkGw4XG/7GeazilBk4WzGthPsVF3MwfZ3EuQUv7RqT0b4WPsq9Ns3K0lW7
SdIglfylnPXpFSO4VmI6aF3oHvaIBPbphpn7lXlrP+tt7yaw+/nsigzy+6Spnlu5VQdUYzkVGqFv
6yaaVVg8AvYKohlzkYfsA+SSejbxLLwBxwv5qCUxZ2Pc8qDPBh2qdirIyMLCCnKtnSB1Z4+qis4U
gjWxWE/+J0n7ZlSuZ9pKi6aC1sMt504uI4qQDSvSp4z/HKDGlnr+cBGKQQVLgh2cYvUUAacwJQUP
lB1Pf3AJHK2ntpf3AjlsOXALPuyMwnboh3zE418xaqHdo/h4o8pNjt/Xvcob5xtgmG7XmGWT0WrZ
CFjKVKzZ3Sjax3ZcD+i1NwhgOQpSo1BrcAIiiRGK7AvgVsXaIn8bNQp2fnZm6Jl3UTvCvIRGYebP
YTTOw7G161Gwnk3LCEXQa1mN4VmtdJmEsTctiH95L/8Jlli6LHX8qdu8GabIWw6TCA37TMZ0rjjL
vzOTmBhb5fsLHPcdRGtjTP+bveQCMk+zYOtCP6lzFapqkyb7CAC5kygiieb6TGDCdPbn2L0/VIw+
QMOe5eV+9TMUEJS4tXliXr4W0f8VzludwcFHPEvEgc/mY3/cRpLgRT4IuNs08cJ4+Jy1l/ed0wXl
Wl42jxFEsILHCX+BxDAHMbmAMms5vhPDDzbOiZURkZ1Hb9dZ/bNoIzvQz2ekKtEZjNfIxvhNr1Il
8y0ZH6wPEAaNcAu75brzBju/AVNO8ojfDdOesHYeqY/mJbAJX3C3sq9akc9KJHVVuxRY9c2DMDCx
iRVBv/FYhJA3GS3p3/rTukckswM9npinUBaCcnj1GgO6ROgB1Mnpxk2kRfRUjb9YUJlKTZlc708b
kk5HM9Lt747GTQEf/2InSrZO3O4VikLyB4jr6ObfPN9jagmt4YbrMCcl71JIKlJqQlc7bHTqPM6N
7u5mNDf+9AHlZH+W7bDU8sL7o54KoZSqoU5AYEM69VHcQ4poZzvK9JZYnxkxhG/I4h0UGepyJcKz
piwENR0EzNWO8OpYKulrQNXza5Q8dQIWC7t9kdbPba7WFPU/0ieQHhE8/sWGdYIhuqzg5p31kuig
pd+kdY82SRx/aaYOH0Bqj1LZEnL8vRHMH8H/bWbZONZNKeP8WBtQ6J9JSxO21HHbOCGluIiFw3GR
rPmW85vgo9HUO1SG3ckZmqxviES69gvkJHAOjIJ5Lo9fwHJAY7opHI4Ie6VoVZW60h2Dje4tat2G
4ssp2+6b4OEB2DafsXv6l2ZmZffTiPDaESUoRyXKvIduLiuvcQnCqQrhG/Q82DG4j4AmSCMjPfmK
kT1mpIxx1l3PjasPzHTsFRvmXCs1qYuaU5NN5qMcn8dRA5zN4QwzgQUuRyQG75Tj8aAlvTt9ZEzA
+7YWjqgFjveQFlX9otlvgnOT+qFdsJ4ky+XVOYgmT6NTb034xSP7BkGgd6yQ9qWHYoIv7GTn+9sa
xaWWs4ygcauJQ08OyWBXrICbAE2nomezyKYbYg/ojfAbrf5/z6rbdMZaMvxZiu35wiQthEqnkGLi
yrl+pMh07e4OL5rrFwpjF3Iqa8RnKzQRQ0hKo//bndVdoUP1hqQooouT/w5z3jMRF/u3Z8Elsq6n
uP+3ULqlZ2aSb7qVt/rnHn90v+Pu8tk5hd/EN1Lq+pZLlBo1tq1UwcvSEhlsAd//RZwiR7WqVkoA
Uew4os9T4Kyf0Q4m4V4zq/ZklFo3Qrc4S12OiPhdEGFh7kFG8zCo3Tc03dLSduT5QxwjxQPWhwr1
/pwsSaGdgqIJzKCcTrFBJTP3/q6fnrIf9UQ6SQcvRyOVfQagrpw2e2cnRC0tSv2OB6q9mbGgHlIE
AuIdG17jsRavMyA4CKwOBRFu8RiMpY02NxpIV9Y+TJZkvS+mQieBRVwyzqaNAA96/e3KkelM7lf2
DzKreVLq9mrfgcSbv477Xi4mlvqj8GdVuGCx6+VkrJyEtnEGSrCN8s8dIH1GITK2qKOjj05qV4BX
YeoqwkCpzSBO1r/HagNcPnI5W5fSddF134CiwgsfkgSqmZqQN2QaJ5pwLF2lmbxBhH0ebFVHa46K
bGPJq1IIgcmU92hsCOHU1V0bSQoPHR7Lvj2WW0Gr86lrCM+rlDGuzQ7O46O1Lfd+OUw3ywAQjSxw
QH61n8W+Y9jpxeH5/gJlyWR+Q2sLAMRVlCBnolBzMqTZy9GmuIQ9PCEgsaPAclCKGEcgSkOyO8ox
n0vklDwyVj77llqr+QxisRZy+dGs4ShhUYVfW/j4jX38PVpuKtev3hYGRJcSeOb2cKbKA/G/80Zs
5/8S8QfyhJOiTIu+jjuqwZWM+6a9Kq/g9rbTQHDSS9avWbXHLEq1U2PumnRXnD4b3ekGypATREA2
maTX0czcG8btwN8vzBwFWjQYMpO0m2nj6HKCssfHlL3PAIBJeOslxgN+farfwwxKH6xe6fTVJnL3
YzrnjXdvNIR86PaL81J9YpNo3yXp2vIPegxdopt68YxS+Ua5Jt6b4B3w9fmb7ixAJ4sEvUOiNL5m
Zt4hGIg9WSsF6Pcm5QfzYf3jmxAhyEt3j2/X+YWdPUJ2rdwQ7uo4znubsbbGL9yviDb+ZSECaq5A
pGUDh4IFubFk23NtK53ltw3YQoEfu/90ha2ZASEoI/lQCuHSR+88l9GgR5HvJnY0B9HiuEJ0QXMb
dhtBSB2iDS6PQxwLbOuaRZbg1tGesq0ZqR6FVneNXJHGxxJncjS2mILwMU0SL8a8NXod7OD/6Y4k
M2fZNrhzXMINpqO8xC+TTISUshpayGiYjS713eNGKcPnfWamzsaszm1HKMK7xo6aOJ6H3/cfD127
Z6lfR49h3nwpI5Tddg/GTLDfvCmHlbQ6KrNmEJDG1G21pyPpX5Zie7eGGgZaA87uDRUKbNCleaE2
dCAYpA/iDzUjJQ5Q5HB633x1wPn9KpXw0r252tIQqXU6Q5gKXE3USJpmfaUWibvOk0YvmmWt3Bo4
xMFWtUdbst5Cc+yXHvy/7GReu+dETyuzVDo2s3ZAqm2mGK8e1dINBulHmE/rymSRqSqeeP9iZcRw
1Ttt5bhiYllLK1ke+0ivXiaWrClJo9o3Uw6dsYAmSxJytshMoeyNcsBGDYhGOaVR3g/bc0RYjllS
/S7HM/yz9SNGYn1+n6ApHKUIVuwNCJdSZY6Ws8kfkU7273AiEGPmIVZ2/YDfjiFfM2Cgj+GLe26n
l8YdblAnpulXowLC0qbZMpQMZ9hQYKfXcUce/OO4xM0kCDrhws7qrLPzPiZypWfCqUXhj+OKPQXk
i+IsdAAGBOp1d8aBGlBrWRq9A5gl9lQEz2obE6ldTEDM+1ktwvWhobvnbBpF7r/0SNQMDRRnHIpk
TGj/PkJS/kvb4pjvBkyQbZzrwAFogOKT65WUbZUXeLeTFM5fgrqGcOjKqM+oQhhk4UhPQ+tTv/Uu
DxWl+TrHMgwi8MWCtSNZJ5sUB6h7mVkYKexcD7E1h8b9quWujf94e7LWFOrdGxfZ3fet9KT/D/gO
ue0G0MFjC4H724hOx+tZfbStP+Lv6yUglm46Y0JhwO+ktLLfoyGgtIYAt7lJD8cz0s9VzLsqg8yF
ZV5t3YEPoLq/ZiQa9+DCa7JqtycWiiz/lCYkcizz7j9pDvNoayhGPiX/iz/FoO5GhbUAqJYkYeTM
QD9hLCqixt2fxol76t7p33SABkf9RkETtX3T8g7aJXcHti3MGlHCXWwX2c7zRvRLgRFsiyrMU1h8
nXlN7lkBRLNrTKSYiZu/DwWMKKu7WuAZuWVRrzAgDGSSBZADyTSb1dbnKh3jybJllwAZsOSWOESf
IhyI9/NVtWiNUSOsLcsYbKxdWwXWFFIxT/MEsVu39FuQy5QwR/ipqhqmXEQycqriDgO3qO8yIa8/
1VCShP7rK8SKwJ2Oyn4bd9c7PSYE/D/OfsNb3TX42VNxX5nfzZgKb0OwDznDIX+UkXqavWYqGKYy
bhpO7zurG8sFJre5aWtg29NOYekXFnihqxGv7w6D8fkY6wSEB86lP/y5pbgmAadK3TtlTAAlM040
maWKN67Aa3Tb7GzB8ClgnxB/ednsm8bkw5D+krkfiHLM2sjnJqiOS4ZF3IaGVFBjT/XqE0hx0+qV
BhqW8TUq6KyypH2Lxg0w8cuFLjE10F9Cnke1365KoEyujE2Es7le0SAZP9GUV9vWhAxJJkAI1M2K
7t90OSRZP0vdMtjp4XBI9K+qjYcJly9mJbiJmQbS4mhIna0Bg/H0aPZqtBDG8oBq7vPv9GyqVrpL
3YYNPlP05J/I4Fyo6DEeUcIalSgVCAPW8eSP2Xwv6NPG/0sVwgSqdEiogtIGGy7b4xLugCt1L4Jz
HvPykLlalH/mSEuR2WQg4v4bL/gvIhZu8Sd18M5YvekyXX5yy8LyQT4MlzpIHZTW2XXYUrgaIpoE
i1hXIcJXnNynsn5ON1qe/SOedqSypXFHi2s20MeNbfHc4919W306woXYstwb7jwFroINxE8aNffG
Deh8IW49ivdaQ5yrsbt4PTQ6WoOJmNuVSEyYyzeIHmAMIV7v+wGjznsXmJ/h3Mxo6FxDlHFoMrSP
PDunyTlmHvZe8YB8tdE3ifD5jNVpFEfqOdjzAVjyEPnRDTlxqrb0zSXXQ99eGS3pZ7XglSao4rBN
IMTSE74FuL8eAwveXyMe0tvSe69YDlERggNdSTUD9isFN/4fuvVEw3AshnMHSY/TyzCxMwyb/clI
OcOwNfZn/5G/wWcAPvrhew0q6XzFXs6JAHGDagjAlCrkYgQTNVYuyaz91Esm0bC33riFwr1LauRw
k0uryHrVdPsP6trljF/8Xg+om17nni6lHA8G9zE3mgicqhM9uJ/r8nG7LqydGrlnAdhZJTIDWpYc
XErDko+3KsQoL7WNzkMoeb41aMEzZBb0gE6uBkfVLraOnI2EfwV7NhMK2qrWkX6GaD9JNJeLqJeY
u8y/5pSMO036Tbxcd8MswMpqA3cuLesv8WT4vyDR2S+6RW5rE02191Wx2IEWoC3DgrfpGwFeP+N8
7yC4VibpummyH9nKjoOjQqL59/Ykz/fCsUAiPvv/5ugfTSBJtK/4/582WDGVqe8+w5nTSLMYfyeZ
YVkjPyq8cOY/k52prQWKU2wQzH4wsFESxs6iWBMGY2VqMWKmeb6R+3chRsHa8z05W6zUcz976QTf
J0ofSuf+YSBBKDgo6JH22OKlmj5DRbzGrNqDO7wZx4VxBWRSQVCVXQenSM9o0swE/wBz/zausz7l
skTuS1PJC3zCh9CYZ/VNx74VaJ61nBAVmdLhM5ncJAQsFam+mYQngAe2rUkcwdF+cP+fCehVsOA2
bLkhM2eo7PpfZG1r7rNAhHZ4VoOcNPBuAwZqkskAHsfGPc8FQE9gHOKDNc0wkhI6eoykbi8voV4B
2rLM53r/mSoNjV9im0znrNjA/Cf9QJyesYHATMvJD18ymZUpwOu2ey2y20dDFrJLA8WwKPo3gBxC
yB480fVY6h68E6hdfAS3rHIgM5xJ4d5hE6xTO5QUYdxPqs4UQvv8XaZN/dhKJvzo2aMhXPOX09+G
ycpbWPHhGNA6739sMbewPR879PWDr9JT+kxkT6l9E73BEgCz06TPLxbST/KZgeuPiTFVaWWN0knD
MyWQ/5gY4PJiRZGdWe4bknxehvaWvlo1cCOMDzYGh2vlam6nQfhtzYDkJkhnBKUVwvYwBabwNX+Q
DNpX9dzuInWoKRRXPdEXZY9yGBvYA7u/2myzWpc0lhDeR+CcCS1yy9k2f+VMaXiPv6jp7HIVCruQ
7/uZUroog3w5jwpNOctKr1l1endL30FepgQYpOS6CaXTCnnu7A8EWs+9CFOi5CpPkQjDhFVo/sPq
T8Qr3rsQUBGVjZyxg6C7Cx0jAzXwNwgMHZbclmFxcnY3s2zIS0qVfqbne3rjPsruI7h0tds+fNsq
ooTlIoNk5A2uPno+DWbmy+X+TmVO269XnCGXXYW0k8BgDVI3uZjdmGTxqboqbqQBfhcKDv6cm28u
nTB0+HAt87fEDC5GpvaSdCr3oyEtKihi3b4OB62mOV1cLFYeCXyKGUaiwsk2Ct/2lWGT9d6M7BC6
2+fh2mSaYcv5DTaDhonsjWIthZVDMSJNa4I3tMmWqQN71Q2wGipISHSaGEmOVDgBhOPehMdvQAya
9UYCwTKRi+gRl8GjbzpkpN3ffKRJHyxKWRvKR3B3wPnAaYeglaVQzBEqLAK8YjQOqrwjHTDjgfoj
O6CLFCDoDA4E31MGMnzVMHLjsit2wa8f7/FGr9b7Eqcjx0Jl3g0l7MbqYAnKV0kok1W4jZK858oY
IanFOZdwBuP2XrsjaHel4mjs/V0R1StcbgVSYooSYnUXxlVDHJU23Xm+HOtfA+3PqT29A8JnBman
7w5SUn8O5HM9AZmOLjlOqNWRY3anxT76XhM+RJO9xVR7aRR8PmhOACuTmoJAWP12TQ+5tlwcmkPj
joecg98Lf0sW+KW8GVITlEnjlQUP8IWu5rc07Ods6IrLBWNUVpInzFOelPF6k/YrZyIC2b6hksS+
F1yZQD8IezVMiW33DGr+haAaavnOfFHKBt/q1svtBiWgk0YeNuuLVUK+GVDFFp5qlzakDxeNRZKu
7qpYMLMtOrK4qz5wgBFYhaDMaXOoX9iqVtYDX5MG+1Z4vY1uVzDKA9rNTIxdayrwV5nbUIkDTypO
dEWz1Ocxa/w1TFbLhtGKMzpETgJ9lJwwhcflg7umJS4FnyEBugQ0JzavqJg3n0ZQDhDOTTTmnEtY
GVi3sVS24xYgC+fB3bcRKtS1VLZpCE7MgGDxzoawbdZ3b3r+Tcpy44rzWE0PnThoUfvx+7b2DtZT
R+U4luTLCWb7v4LSKHd0fuzBD+cRtJW2vTcAjxqgUjJnKdRyhl4hnHJddOFcZVJUmWHj4AqLo7Yq
t4wUcVnVQ7RY6VlGpyUSx2MPaEt1voOSbjpSjd2qXNVQVtsEDc+GDS1SLeWmFGXN12tEBM9fr0d4
PN2KtwIbH+Ua6aQq8O+B18jJfrR3yyjo/lLDC6OK+wb6+fEoM28MRyYi6dKpWpyUj0XKzWCgTZV/
4b8yYxQWMwKCnS2EChdYNzk8FNqmuaoExz3pZ2/M5NT9vYUUaBrWk6tXAaQR5pDWFporRP3YKFHd
IT43M83TjaK1zptVKl1DIygWBUB7MjrFqZhwbx6xU73TSjpsEX8RFr1mlmXM8lE0lBFR54wj3DxV
6obcSnyQtW7vKByS/OLHMv7gnXgvkwgJ7DXs6x2Nz3devFSrZeFFsXaqQqHYum2VhG8kkRA+YUE/
ngLaNwuBKDznK7hAJZOSJ5HvwHTldLwY3ges+Wp/0/Z8KsLMOYJIY++kNgS8QIDJofwnOeouSyXd
4pcnJuyrRlGF4o2f+J9clhdONtqhAO7xFpsgNZ4wRBw2ovn4Pc03qq8vJP8n6iBPtGML+uEXdaTb
Pgtopfz3F7gw7BXg8FUCLb58WJCyAAC2w0rBdFXplckea03YkTgxvYuDyogXr8ZMkZS1tJl+o3do
u5QoRkFTBxS3xC7UXJQ3olZCQMzHgQqI+nvT9T5vOfRkvGDxJaT0W7ljayXTc7ueaXb9ijV2R7+T
tQmmsNx3nRbZd71neSoLNNaAPB9ysUgUl5jzhOpX/wiwsMg94iG0ESjKEfuBFqwOSFY5zhPKRXoU
2j1SzI09aEkFI2P2SYS5bjjCuLofQoOY55S6EuhguIcKpMft7zNFmS07NuhG8fXOyj9IWqrkn64S
bSlfJNFXv4ArLt5nuO2bt+AKMRE6dS8HVDIBO2m1iL5/OIDNCOeVI6Adioy9dO3sKGuOV9whXW1F
oMBKwmvVAp/q9tyJrj55ejt/ja5D+WFZbA4adX6kvDux+tALnua2C5AxlwraOiWoyVZmbOM2jltw
W+PBQuMTmJOwiF62ItlmTBRCUHQlGRyQ97FtMoehNU+RsDIJF5bH9GNcat/iwDuzvdH8zaHMqXRI
E/CTM7avFrRqpxLG/tLaaW0F3VoFntwCENCSp252PtyYWNGVsxWD3guVgY9sl1U1dLsepp/UdH9v
WSZq5b/0CfYQvaK44mJOzg/J34Oj/aA9veLtw6vp/DPQHtLGNSOJAdXiNKkt2hSsf3+TQQPhEE2+
AfINOwjr0q8edb0XhrtS894X+FneUv5a7q6LNhlMm9hPXEDvd0i4dot47+Y8P9Sei7h69Eao8FGc
VqitQpyGmMIrbqhX7AcY1bwmRLdV/P8NzWsx7aVJm/1Ch9oNGav7kwTfVK5XOo8/Zg82Seak5qfY
ImEFlVgvhh7gmQZPFhEpfjg6UQWaMt5IBg8AX7MvAyv8KVy70DyKqOPy1Lol0/SxJoByX7bkKNAG
CKVpiXKiwWIyikbXGaBo+T0IJT9MgByES+lUDJxzTuZA1elTYilYSqWMMjUp8JA16d+vgKGpqcyr
1w78fNakD950w+Kd9DSIWjs346peLS28yekbkopR2J2M/Egac/hPkbOj1FMOJjl3d/DSRFaMJ6kr
WZsQju89IV2ak36Xu7cVPaDL+QthXWIhStQMYcm1k9ZakGuVJBTfKv9iQzoEV5jRtgv0F/xvOXV+
ybMR9R9haD9Y8zSR1MoTMR1yweSivF2Ia3MVaESwX6TcgvILXMVUIQNexyCylR4DCOlyD2CsTGtg
OYCwRE5m8zJSV5KhWY3bqe/DpHro7A/kvxRfdi1co0B9jSMqr2jSus1POhSDksaeCrTkAI7vvkut
AmuJgzpNL+bcfZUKB6DDEzp1pqSMn6H2mLXz7rtWRchH9yJdmiJqWT7U9/XgUe2QMtFri21uPdOn
43upSOEHxMzHNVJ7OQQVnk0ZQ00sekLxlEq2qK2kxtOdtPzeyQ930wpXD+SDFHJKZ0LOnDoD+PKU
JuiFPpRwqhMeW6KM2hpRAczzfvdejY/TXrK3U5fhBwL8viFxsDN8AugmfDAnOg/wA3n4ZGPD1Es3
ImyF8zlFNSnOng/WZF3E4rOAE4kkndC3tsLHLNWNQNo3rxtkoWhOvHTQ+XAFEagH5Y8700mr2VFL
2lGlNQFId/lMKSme6Do8gOrIk6l2WcloHkOJFYZWK28G+RW/dEewGS2K48SfSeH79U7FJRAwDCRp
P2dvts49c0xsUBeieaGczLcwPbESiSupMAL6QKxm3ZIkRujSjGkC3ZHzGuLQ79eBt7YgnmzNO0Fm
Jz1xUexQWqDx0RKKWBFnoIYrFP0ja1r87ymA9oYvxyIlzvN81/mYGv1kCNbCb5QvfvZXdPkXURB5
LVB8YTSBDCHRakNrMVkQhi3XRa/0uhyyMBWD2N95yOEXRKLxlxVvDVjuH8nhaTwZvwfR9mRsHdR6
LAUjFLD3xz2O3OgpSCtFJLuoITEsy0dm7YK/2sioCF4OQwSSiji0x8Ki2/nPUSNJyUv7pAaHgttH
K4smDSSlUNNieiNEw3MY/Y2o16q3eERQUeIvIBBxmVLFpiQS5pqNex7GVWzyRzczwkuqj0Ikinfe
MDv6BEANlG10U0ORkXradzh/co/sx2C6Axg3ydrueoWSSim2LJJVwJa8I1CwH18/oIPtbCCkB6qR
HBNu1fDQxXoGZJD/4F18vJTkML1m+2eQhEHB2CYLs5dl8xilyop2ZukruM5XKxdPzPmYauIJFuvH
gmf5Yd4jpDutFRJ0vpkjXr2o0FkQIp9RXL7WkNNT6qMuSy6A7auqNJYlCG2sZ0ULMCwd1NMDFREJ
i+EBFpJ5PGJx6Yirc0i0aIMsb9YfjcI3VY6xVYknAsFkL64PS470CQsXuNji6AG1QeTif30zs/GT
Cm4FsjCcSX+46QofSS7PqhUxlpU1c1BnhDmTeKG8fvMyELtR7BleXbquAfSy0ztXQNbju3242Ll8
pnbzg5pBsB5HukMtgaMP5Okey40CDY71KBAMScwM/fMGQZvmXf+EgDitJ//P1j5we6HxK22Jtoiu
4vzAR7dfypWzKog9XJ0Av8nfojxSmfqDyB/2L9QxMmuoO6GJ0z1L9hNE8GQ+6lPHJ+/X6s0RQ5ol
XrF3YFQyNywoxEp4PSXMaUyBkCXEQsEJo9L+em0bXZMwK2DJdl8wPcHl+AQDeaAjHLgSSMZUII2H
HHlmoJ7xG/ybzFWc1werQRA/7TQXPbFrf1gXPFf7Ii70MvebrBlH7e143mbVtjgB2KORTxaxP+tW
Ke0+Sw1SU4G9YwMotCyML1c3VW4c5wYyeE5tob/H4n9lO9PkQIpTzIbdv2RUC3KCigkberSwTRtG
+r4wJhsGu2YR0kCEu7mgTrET/j6NEY+idZGsKH8eWvHEvaYhwOYHq3gIv5g4dYEoyE6T3SJhfLMA
r7UGcqsQxDLv+bwuV+wHDqAHnT6d4eemskhU/xdHxkAJ0OWxKNv4nTI1r2YzWIr45JO14U73c2mq
Arq7VU4mhi85nFaJcCw/Rs5Tt0OcL/9Z6FBg1xVjMZVTA1xfNrmAvXJXwXuMgmN9zQokbpAUVQ5n
DvFUlYx+3YC5gX/X76iYIYAOh4spxoSWY7OTmfkoqFaxs9aJ52PEUAFAqOQ7J4lAyrs/9QZtzfZa
3qQvfxHzhDDnqa3wGPw/oodybU/mgMZNFL50xdEb2lt+8wFDDzJiuEVpnYXW3iUM8rnWbdQ6goLv
dxaL/YlmD7LA/55xVTx/fSzqsRR9yKrnTF9Jue2LZdqn9M1rHmaB/ljX8Ksd0VvD5LJkvutSqdaC
OrX774hzMdZDC6OK0SmMT5ofY68g39kY8YKHgxA9j1M1ujMdCo+QjOcrpaPUNxbMWwf1Br/ejipL
1G7Cr1Wxl13agORuW1OfE1rqUv8qpSu6cRj3Es7VEZ7BdfO9zYqYlLMiqb35jHTx6BGgZ88segJF
FMfdC3ECN94GSodj1jUGPI7UjhPnqJzHHQU2QYFrWBPScS3B5LjMON7IdFHHCS68BjD++bUu1jNY
uKKVoMpNJIyMQHpkFG6p96VVb2aymYphs3l37ji6hNKjiCIu9s1VZiygGFzEGx7Dz6Ajs4OVE6Jn
hhT1ycElHd3mY+0vv9LlcIwxGpdUWK0BQBaPdfVprgxq+gxPobwTYUw+Msp/EWKlsMOccpLlr0eU
5s5/ZnvQl2uwkMeOUw1wYKFHFdmdNS4rwJm5/0XdzQM2o8OLKoaBxhmX+eiw37wPTS/yW5VbowBw
rf5hVLr/JVthXnzzojyqjcqBQ+AXJjKhZclXvQFAHdmoiiBGD7aZoZS0kpXlOBMkRLdSMjuezejO
GAJcznaeTWUE+g+qyIpzJG2o9o+58Ug3O5D5QUkrXZe8JTzg92nc1wX26vhbRcABuaAKo7uyc004
nfDTc5BIJV9PsSv7ci6rLLTc02j+hHFkziWIKfKzLXpVd99UK3qgMq4sWi76ZUG/33cHA9W4lZN6
YzTFhriI0c5VR2VBkmVGRqr5/n5TV7Vbd2ma06fclCB5QplCaguic6LOx6/RNRcldA5XDppQzJ6Y
OH95EsperROQ4BhfXWhlYxPtdL27C9CRCAjJq/gZlXA+5bmltsBdc1RFY0qr8BjlXGWnqkwd0+Jb
mrUzMI0lEPtZVxq6no638jnsG5SCAEm2o3n9KaJFcYWxcZSCCO+IOuFpHYKbirhaQl2usHHd79Ok
ZLRt7XOWtfP719AIAWQK4A0jB47IeuTSltvZRyIGK7OUWKAX6f3ShsD2fQR8vWN/J2BljWSLzA2n
cVmR64ejoojzK7Z5Je923Ch5oh7LL5YmWP0pJzWo5NpNwztAFwJDQ42HYNq+3pLlSi7sZQK4NleN
YbEEvEEDcgeBK1eBowW6041bCJEnXl8nRmjyhAtPg6SnJLxy5q/5EpbnDQ/CH/CRytjr6JoiOi01
v4M3u6e+j5Q8wIUFMHJP0tSupAArbV1UKCmLkm7knQeEUK8uULhQRqlIZpWehdOq7NJhGfGTAqMG
+O1z1d/CstX4B8FTEunIjyaZT8mhcx8iOoMg1CM4BtdDELGA7TDGKvgS9Yn8yCw+MMAMwDntdn3u
IZNNRgfI3oA31CVkBy4jyr5baoU2tk7u8Nibo2Nr8DF4Qu15oznG0Q5hpZUmmfDPnOyN+818mdIJ
jBr5lniCXbiR7VjG9dSOZoTsdbcwXBT/f0cM4nM8zLLlC0xalRGRg2W/2mjXCLN1DJ/MId7Mdlah
BnksZe9zWGBvsVkr/zBxns6fjoX/prKLvEBpsPGWGlMj0fFbfQwX1qRjjJatxpXZ4EE17ggJKNhG
ca5EW6ymcOvhZKB0jTIRhkhsSZl/N32A7NOCiV4Oo1VaYLNq72SM6aAYbPgGG6yu5ME8MyTwK9lb
8iPf/aJ11A0GS8kXecrJpZ22molfW4Reh45LET6rYOrMm07YsWcSnO74Nz54DTt7L/P0FoXF+e94
MorFI8rc3gSF4wLIEbREHMTf7r1AjVDRGXihfNaD6i2HB1Yevm1VmzCAZj/zVMSHOmHTu4zgD07x
DzghpPE2IjN2ufTZn9KSGWQPGC8Mr9LLwAj12cqoOKGcnOW3tu6yDyc7+VZdrN2R9GPir3r9giR5
cmfaiMGqPSffST5yK6z7IpzcJt8wlhayVlBhk6zYBMLyVxieTqOpzdLcB5gHmtLiPxX53lH3t4Qe
Axb8Mbk2B5KJozJQ22G+Iu7px2ebPDO0NP5vfkfJFpo4xd/6jDCE04llq+LHs2qODCYn0AhO/KMf
lKb0Caz5Ts9k90bc1vYlfl0NYDABqWafkbNJP7Tka2fp/mS4xKrZ2HQGINr4snDs4M+tywr2pml1
Wq3Jb4NrDsFqWjE6peQXQMrHc58BURE+YYZNTEdTMI9zEf4GwtQZaZz3cu/K2HIuc09sXS7W7zsq
RWYHEuVZByRSpiysl7BAD7wlIV7+IjmxjZxkQepPRCZhtt4Mjb1dTENpQYFKph7sa7NUTqwEhuWd
mnjoas5V+xts7GgtBATtarFcBhQHnTnDwqcUELvNtOqKnzqE9TrewtlsrE74XcCgxzSs6rDwFEVD
TK68d33J4ykhxV1gQC5I30Z7emuYW6Drhgnue6eQoTp0k5UAcbh3+dX4h+ZDFaDaDS6npEoqwDE1
em4w10z33P2pfGzBu096ULuXGVBM+HqvGC/1MYUi5PGMipyUwUlvILNd6F58khVqIst4IZqEyFeA
lee+FIJAWONCZ8R4CJYfIpsAUf1jIUA32yDCbnLPGb/0/nFwAaBoQ0toI2pN2huMIbgfNFp/NiUd
UlmamHS3RzR5TVpEw5BzqCvTcPEAy2PkHnEtCViaAPWyzh7L90QCHe+ZJuYNUhMmAOCBdFGKb4Gu
WJ0VmqnkcPrl1enpGB6KqP05KrnsQCyp1+/2nMzs2MUa0+9YjzZUPyJO0m2bMYHtWwF8DJTFEY0O
bc+n2f+hVBhmltOqoftHlPv7R5oZ11IptsJcOKfF96OOQwh6BhrMmHN0iXcXCTifGBvtk/Mm43Kx
fs0tW+Q/S1ImxQJV7xK3AotaZD7q2Or5NHXmmKFldYkP+MwF7CGI1UOMGYe5PydbHK4lGCMq0J3f
9W5YvyUZGmLZRxWtharTbPoRHeDVcq3zdhObC64dO4mSw+zvospg68ogJ5Ys05SZ6WOit7WheUn0
a8dI0B7LQlOJhnbgPDgHgk+UlisvDZtLRjgWGKIzJdysS8O5ifzMEqtN4Kr9+PYxxPbx7i+JN3q9
REAA051NWjAs2+vrGm090UYK+VqH7gQwS7w0FGiFVyWSmFWmEBXB293r85vtIIh+ZXVxDthLYllt
ZBTDErcnNEwjUbQb1FoS71NpXB3D8ZIOLCkL62QIIRrJcMF9/fROxlMXHgGO6W8Z/AtGRIChPV0j
ZqXj7DebVTs5POl1RYHXI4hpZLUhNlBbolmSBePred+9VqIHX5hZ80Z8IOfH/m5QH7TSRUoPpJqE
dOdZPQku9GomVKKJXob7IwNG2PoXdQiQ0+SpTpM58fLBHJSReDXLwjhJi8A1ru7NuqTizGzCF/Cq
Hhq8sJ/sn/kE9QFVk4unbGlRTqKrxzNt9BZlAg96+WoTWuxJnb1ICMeMNbTfuNOeEH0HiPS4DXyl
hO3KKu42pRAHthZEoxhpepzegohtuCmBLCG7/TbVGlgnI9aoxOK2X78IfpSVXxHvHiPc4nsrPYlP
EI/yFvUfh2Kw3OS/VDNrgrOjSbff8lAZcJU9K0GbMeQW+AFlDo3PJI37n9oi5pZosRYW+MzorYqS
oYQhmVRmtcpoNxUJu+H6j28S9xvZ+SMaxYkU/OBmE5klGNpNMDdajsZsSj77EyqJnUc4WbK93G42
Y4+xMVVd7+AAQoTpCwXVkk2XMTHjRSIZ2kOSKlzQ1wu+k5xtsCPxDzIoJGGbv7y8t1t2WsBuGRU0
P1oh2UG+YiAHQFA3lIpgbdF21X38moeMmN2v1tBiz3wcGgQxNkOd5f1vjcFnQOE28zIQSorwv7pj
eQsVMF/OJ/+yOfmdyXYun2Tiy/cCZ8RvvaUra3Rp1Q4M8iGe9HOObvZlQhL+cYVjAritNIMT2Ypb
kuFTRDpTqfkT+rUzPkLVSiDzIn9lIMDaCGUb5YeMFDT8918IEfvQ61cAK3aMzlRUgEbjh0rAAqxw
Fet02kg894WiBrqBgXWesbaLHR6oGKlgRm50s6aJbfGtJ+IlUT53cT7fy6hYyQicOyc4xdJ/IstT
i/F5Ay4g1yXZNBIKmFXhDfWVjq4UrjBI6o94YKJ7EF2SMiL+P7T/45Dar8on9AqqK0Q5xD9d0vNA
/KL1+OSf+nIhCZLiEZUqxMiAPwvD1UwbZG6vHybkYv+1umnSv8+47rqlmgOOOIy2twhZahj/PPvc
TKztPdogJI/2Rg2Bdw7vbvmEN8cOabzDk5eCxsHBK03N3mBKRhk53Ec0Y3IoOfPuD7BdqnkIDRLZ
fZ1ByvSDG4WCZwMYuwvX8varCVonx6E8KtaGh5FPQ9whirhfZWFta81Jr20cG/0DbICAqFgCRLPA
+QvNZfdQqTqabGTJtjtHfOLTJ1FL/kCCFRtcXfLJPuguT63uPrb9FSHII5JugdOiF0+wn5aVOZG1
qegqLw8tp6u+BKlh4uBdu2EZLKUIx7707YYRNoGvD/vJ/akOKziCzoXWYVUzJEOxUY6CKnr/09NM
FnepbCzC0ez2WZrbdE01xTbBYYdgzv/wKSuj2bKjAK2tn5JaZxlsTqcSbddZr0Ao08oX7xSfSYsO
+HdZnw2aR8dedCKXtr6Xogcedcv177UKUdGrabgHr0GDTN8LtAP5+nirjrL8n/crh2t44RGcyh9X
DcIXGditc/CwyxP+8Bm0N7Sge79IRFiq4opVyI/tObROpwKHxXlV6n7ItDITRqkPU+9YnnEbZixU
6NAuH4JlSprpuSNxqCb/QZ04th4FT+nbEU3ZqvcVWRZYPywz0kO0HaQ2YssBCoqWRb4DUp/wrx1g
nlKHi6m5ufS63isibsql0efJhMR1p/TdSMRlR0rCkn8AcpRMYYzBzT/SAuyA9Zp4BGNbcFe09DyK
Tg28rYNi1qWkKiuZbPpDscUKUUXRUryZ36AaZd8uUYq/zyWdlbw+wE/M86UIkcZZfxkGGfuHHE1o
vkiorjkXmXIoEOUzCwbXp/IJjEGCJPsuYgffJfHkidfB+PvHZTArQH/DdhHL+9n4mxofw6dR0d56
2VH8rynDfbO0HO7OHXVMNJSin6KW8h+AOzddNk1Xl5UhjUQCHI/bx4drjfza+lVBQlArGen/8Rvg
ESt9qeOpDTEfJTUsBRxAtXp2H1CV9fbDQdWwadnWUuHKUWSOXguQy/CcaSCOdsiZRa0YYwa9bgH+
Zky4HYa9U2LyZq+G/PhdWNpuKjhQ2F9nd6hBEBXaCpkbY0ZEwSaxjo/Cv0EXzQ2G+hXAnSUvFRAJ
bTl08mlxsTxaiAGmFQ8E1IGGJqXlIX4wdn4yw6hn3wdFadI5dCIngF4QWqNsVlmpMSAypE3aHhBL
73mPsZHvU/L+tCDbRK9R3Vk87SE1xI3Sl3ImNW1WxHa4ehF4+ToYQyo81R3oPFsxNEulrXo5luah
DwlKzHCHERjtK64tNXWCncdR5OyyPbev5PHYM4rVev0Q/C1RccfdH5sL92e/iv60f/Yl6JfIzKo1
1ieioQ4BVYZc22Ud5ufillR6JzTKruOsHSaa4p7zbyrfOPz+OFgBnBmjPG3OzMokY24nXNzctdm0
3mCvyQ+lcOWQKKEvoIh4WAZGJNzOQwu4woEoVVO9OvBV+nl6Kh6VxE2myNKltQmaGXPD50zOwrLm
xAS0NhURH41Hb69pwUNu/Mhue9/Fjse4Exk/EZHEvhJOZvEK96w6O9CL2hF188dlRRIhL0P4AEbx
4Px2D4BxCjijImDhWEfzPcWd/XMhVRz2xEOsjb1APJqouK2W1lN9kX/cQbICx4zK34p4fJ+egRDD
Dxkp3KGIqBVG6ThTMzkqb8i23uXkISHh3XvIha72VcV9MfZSoqzIjMnk3TasgSZDYC22nGMiV+h6
BSpg8giMApwVEAnYL6YxDWednejt/brwywYwb/6AWwohdLsE/4snllBpZ80rtKPoYv6VRigDjgHR
h7CFS/CQS7ss0i54USweZDBdVNFjV8h6nU/v288Z+aBOQZ9ZmHLRS+IP3IO/vPm+f3Sn7x/2Jn5P
nKPKWkQyMuWVlbC9BxqdII1X0jj3RLqzHgjymnBwJ8AL/CNy8d/L4JyBR58zyQksFCjdixJSOqgx
ZrcaiR9XxaEEbSIRUYZb4+wy0jsaBt/U1HosbbaDD8+qbZ1RVUlPZoC3l2b4cg3N2OjYcox1Xtah
a2cCFu8Q74ZVhwpNpdmHBBh4Ri8pT5aJ9z+FawOa4x5WxJzCf+Hpk/Lajid5VaIihuSd4skIHd/7
WFDHjT5iHm45OOTHPu9SRuRhGwde3kN48OpkiQ4OrPl1l/UJNoO7zrq0J6fqG4PsWh1qkp0M8KGe
R/4cmKzgASZmSOWr7oHNUTj/N/DdCVN/cJ0N6xCilLqiKRdKSl2aOEEfzpJRssD6OM/vQnO7XMG/
bvuzEIbbnq/Ri6rEs4tz+I7fOs+lF69NwuWi1DGkIpMbGadFPamxf/agVenDanLV9MsXcFV7m4Lp
hxiP/rSY98aNx/VE7LIek5KmefU1KDvWNRUuy9DHOcHsj9xOMe2YqgJndHsluJpirkaLrGqdlPVN
OBtj+3oHlr7Lergu5NZ74IwatV16pL3Ti0hkvrFSk2LQcctC7flc/TDJrINHhnYv2jj+XiWdBahy
k7O/SJGfVBq5aUoFpWJlkt+rCxARYhrFqNVR8dI7MHKeZsaIeZ2rAaxJf4yq4rEbotwuJsFF2u81
/FDWtXvUPK2aRsd+JszKGD+0CoN7sIWkb1fK2GbPNE/idwoF1fPdwtF/rYJaxZ5Fw4Imedm0t/oz
cgvFCxExJjuZyt8eGMQxWHDpKiarxQeeD+AhLJw6Z3DeGPxBwICVsWtYybAtOWVx2heXB04FQDsZ
5SOgtgwhtcvMKs67RoD337vnA1dMhKuJS+NUYf7erWy5BZUgaialh3IbyUTPKWkg7w3Dbi4xNlb7
HxnwOkuNbLw/KLBRWjctg/R4tB2e/NjFf0Yj7qyc9g682DUcTD3Iued/+RGoP5PYU5ob98rozbFI
MSsmW9/aVKYuioPz57+Xw5QE3g+LziFh4ahNwy2+Fc2akXFsj2/5Z+N/C8lqDoHe2O/kWNhpWV5P
SFd3PX+RzWHuFctojEVBo8iLtqZtddn3hMZP3Hh2YdwXGDxagjd1oiDTwVJQioCKQJM/D1DAWvMJ
dKvMYZhCaAYCO1nWDwnBlvWiWBUnzTA/MxdpphwID4GrITg3v/8Ba/ryRp8mw1eJhopUTt+Y8f0P
30aRFT/FRjmkvG3sjAJ9oi1+6uXjcuqNXAIxtOqAnEV4hmZcQhA17lvcAqpnkCGLtsa605zUEg46
3uy2ZxcCeAFpTIWBGLvFQfvtL9UnBFzg9LLET4efwE+2s5PioDRuf3U3203aKPRv7HuEIKRvAfrm
Nmaucgb2u68C1swDzrr/jbE8KHLsx/a5OfMOB3VHj3nSYqBwfBptXTKg7Qq+4xEAXBe9AjBLL+lY
1K4g3c0WwlaZaNCH6JtYptp+Cyij2yRmk9QC02Xvft/kZmFDg62JtBNUrWjdyguoZ1lobGxbKTUv
MnoO/aUQ7/6WN9x0b4k1ZorqlfNe3np/9WEM3/37TbLVIUfPQJQIEUd8qP7M5IEqLDHJLBp0OFhm
0EmLy76TEBOjr6kPRPPhcmrSCPiedRNQSNzyrogzcuwlB1bp+ET0mwOJwGEdLsYpVl5kOhQ05ohe
Dv+NCtJ6HHj74r5E4uvH6VWB25mC1zlqGshbjNeMBxRsKUom0B9O7BZzMCtG3S9bf/Ojs8b92yQh
KSPibnR065QrEE2pVaUVGtDMpH39z7KkBpQSudXxBl08bUp/ZRnT6jJ0dyFcHWYDw+Y/Rtx1G3iN
8nRSIztYb3Rqinc7sm6Sekp+DmwcmIaSNQ4yNvtPT3/Nb3kQaWFbD0++dWz0BYD7tmaL6j5qd7LF
4m42Q9MYRnFqMBtF2mO94q80B0AIM5kjaflao8Q7K53KWED1sICnqnbSb/zRGukSD2BOQghT/V/f
4/196TwJzRyULSnJMXkp7KnkL/Lh89zA7uYoufjeyPuGUhSw4DFn+U+MqQsWbe3T9PvdAFH5ILp9
f/ImxXYpmr00YsNPHC38zoIjF8GL3DVsMTTpcepALkwOd6Ll3VKcOwcG7LY9cfndIaY+RBoNrVR+
NzQLnSqVXApgHIcD9BnU4La2ZtbT+P0kXrAfNYD36kvN4pRw2nfzacPkY7pwk5sC0JrncVt4MWwQ
YL6Dc4IOv+JAR7D0LGwiChLSt6ZTyod5+FexaeJxpsLWw0Pyv6vHj1tIocSb2aB6OUM1gpoaPdyg
2bYHkgDPE4RuZr2vKDz9kWzHfgKC0XN49exmRuy77v9TlD5QarjzUJWLkBy5bM/1mcs7F0SA3IKR
aV6vPZVs1TuVpJ2otMBA9ocLSb610QaLJEnhgD1InoyfvdmlRBFc31DDMWJxSvN7icSaIkfEXOUd
NHADb6rzgsBdQodNiDAJsPA6Bch8QI/tsaX/6gX2JGGQWr4PwUARppEOEJsNl1yonFq6GMbhQiiC
yBRghyA09IouFXJLLOMAznrhzbO9T2N1E0rUVQnsOj8pXnTmnIJ2y6+rbCX+/o3X7jwMn3qvbI+t
r0hJB2crrwRHU4Zmitfh0EFdtPieFStyzjDRTDdAxHN60RitHyqpXapM6nwWnIxY9SKuZS+KnXB9
9lkDeh8ebcKpO2OBXAgzZ+Nb96dOA9BH0KdGXrpt3to5YgA5urrIR0wuJTD5QRXzcQe40Z3gh6JK
WoW3W3TTXeGHzrI2cGsNAuVk1DFL/yF1tynWNwrJxagLLL71r+6273Vw0wGTTVuARXlj5+aByWKU
tjKltdJAAiy5A9p3ar6XAGcZAmO5/b1De9V74SASq494I70ZpmJ++HQl6r5QVr6f27V36Q73RmVt
qtVNFhhl0uSWE1l978qo+zC8pmZQVJmfrrWlloMAkl9XUel7rHoPQUupvz/rFauS3P1twRZlwiyE
LeECYaUsVTdtD3MuL6Ub+ks3iyDJhlJPLI/UJ7b5Z9EQ7829ByPMhB0Be4z6N8rThtzD62fD5D9a
mcZfk4ogjKSdHfStxKbetpSfWOq/Haf3tf0kQP6cuWtAReYlX2mgITWVWdBBwJczyRfqpiSjJZaq
o8n3hExIwP8iyLrE4UttAhmZwf1911WbXnFV0cEEEqgveF0huyT9Pyadyi40hvvMIZEI4OhjgHd0
hNO9E92GH9oEdXKdxNJJguOIGSEMQWmjIDkJGIZfY059jvLHWl77o1ItaxEKf97oNB0DmgyTD3Bw
IAqXHQgzUYaqb9ZLUPDt8OZ6NOqfiPszVFrRsA9m4GSRfy3YdyxWWJ4KKxfMHY6cTdZcjVvoU/3s
DRdh6rGvM9gizafVGhrHLeV7o42f6tHmiRL4qfMuYjDVSkEROG3qweVTquCw7Yb3nxYeAOWTjS8Q
zfeemdwGRzXSiK1MuIG8ig8vljdH+WkRPm1dLNj9PjnO9Wy//fiW6s66O7nGJXUt/YDkG0pwyU7h
FuQVocFopnP4RSbaRnSFpcp1IF3q3IMsb/p6l9iyqmBpId+AxhOu5MXnvlwcCS/a5fCvgD3Drk9b
InclMnZe2DyUwZ06x8QrVWiiOxVR+y44DHkPdPzDYclQKHSDnUZiLvLvq/tmtVJARw6XGf9vnoaQ
bwlXArSoVAElH8A3B843w4NKJ8Q/HHaz4qaTZDxDAlWX4j0lBqq2USx0rOMgRSyzOJUmSlr1Oger
tksxo7ECz8TSbG3HTNKzPLO2zD4Cn5DW5Xm6/HrsWwznsPDibJ3xdH+q9Swxo4JKWyRI610fBaPF
k+u7zUF4p0RPMzJD+9XgFQbV4iullPA+MkVSBfqAdGg9SCQ00FpR2tuQuCjW5QkxA169BcEHZYRb
z6e0h9G5DLkktK4vWRO9y0FVhSU8f6xnd9udjhTBtHTLwKviufYZSQew1Eowc82lqUffYbOfsLv/
dAq0XnIi8cWe4dovjWRo5dKkUXlC0/c+VuVhoawwg8a391oovpVXWyh75Qjg6PdxvMeXnZsAePdI
s0JRpvgoEdzqQYxvR3l3mhDPy+/iytzEwHFH0cQyhet8WKrcnJPwbsUwS1hOaHVF/w6towbEMjF5
UHqPnY1YC8IWG+kdGDO+kinw36mB/VU/dDqoUeXHJl0Ma9ovm2IhQbspO8pVtbN1cKr7M0i0ajWy
XRCnREekycm2uC66orvInqrULrqFbgvuABsxXh35P9quYjZlOvxbOyAENpNdFKccBqEtp/fulbF5
KCN0o7dykPZNydyoGqcxIF2dYpWjAOBmixDeIjmlMJqBKJ6cgdwaHMRb2dVVS2+MarHuxC0v/DHO
h8zD7mrodqbW+OAHxPF5htePsBgtVlGiduLovKuwQl9vDhBzXSX5QJMxHWL+Zz6ooeBaz4r32QBW
vROl4wKiWGJj3TPc/8ea4FwE3zbv/E30LWbNoBtF8vDhgvlKlNUvl65UfCbvbDQFRt9Bg+yke/XB
FYe7VS3IHI0UpEddTFgxiIXYlVmZ7XlEsW1dG+LVrNcYO83o+q0QnvSXM31wYkzGi2/BEm/Bi5D3
3243MocP4hhbaCqdHvqt2xDIftpGGceVeJk2mOO2T+q2RIpx8rWVCW63in4UzRdzH4yvYOZb1bce
WJtwZqhn4do0ZRaXw6opwwXebawf1ZZoKa3lwNNSZSjKV+qa73zU0MJl8SnQduaaLc8DX+Gc4K8w
EO87k6JDDIQYx5PtIZt94NacTUa2KITb3aMfrRLPuywFsX5caf1no7PuURA9QWvDLGYRLa4RrvJm
XTJcsqtWbnKh8OZYiH2/kUxcyuwffIUPfswn9g6vm8VoiQFb+OJhAOVZaSDwuws+3JSlyMeury0M
zPkuVHR/n+wvvRBbW3m9pmrLZF6w70jsTiAGjl29lX6vYYFT9m9gMjCd9kMhPX2X95nuQN7Vt6w4
kjXMyPK8ID1qtuNQ9QaLA3jXV1rEFbTwo6LE3Q3Ru1vJUr1aeyGN5Pc0m17Q9OHdmF2oCjWGr0zU
fvs/BvEJMzS3ah15FkevjBtd0Jz5jOJK9Q6GqOtrc5lGc8sh6BIs1j6UTZUie2VpY7UhECIGslIl
eSICubWsf/WASk1WxiSFt4gWzhuJmYSuYMN/PnTKvoJNO6Inui8q76VGGRPEdDIYMAg6MJn/1VQT
rDGCOYgIhZkexDRrlKaWzKeDgxH6akQv+3OES1mUmtQl0S15scmlYPvRqrhCzilnB0Ziw1KQFKM1
W+zF8ZC9SDuP7ZPsNnDyK14fS0Q53jmO2Tq3ytPKs1NsyVHhNDMV0FeTrGTRQSt0yUb5JVyAkrhQ
l0n3bwyjUrRaSGuUMr+W8OH5tuTqwLEm8IX0LlfG7jpASbeqLpopN4s3UQKmCBiN4LyGyIOqrkm8
d1QhezcFCSO2wARCbLuuBIz9Ul2CNombLHLvKlj5f970Fgr+0GaNntdXxAouSv7bBeiss1fe2ygX
SZ6dto2Gz8NEB4K29sqLK5O2d/CArCqxy8l7WPxPFleoz0+bFrB02qA6xxvsq3hAiqWjyhBwkfN5
uniO8y8jzKRYSDFCHAlm79y2tNIlwZLyym9mTEzbtzxS0dzdrJ6lVl9tShsdYwLjvH3xA0voMFVh
s2EjYcZaqGae4ppMvByDS0RL9R+i5R54T3J12j/U3xmn3tz66Ipij+DqO5WQFaV2Xjl+xhdwPy5N
bOPrSs1dkkFvloRX1s+d/WppaxcK3SqKdNLMrs4sE1BQy4+sk4fkuvnfnI/Lk6OEXSCdMNSrv4oI
r+UIKQQbeUMNUkvrJZnvRHTKSWpOJIPqtxYWovK8IBgcQM3JcXT/xrVg9GG0uf07szLJwi0oNRVm
Or7dfrW+nEoVLS/1+QL2jMOZ3t0gi0NikT/dq11GWYM498wa2bJDGyytT7jkZIJdrImKQcSmeAzO
dlOojnUVk/ziMxByCR6FMgscGq8xHn0tCxaSebW1G5QJWUJ40ugxDX2tJcrm5gDhX5LfABm70GDg
XdX8tT5NL+lkdeaNvtkyet+19NYpRAbAv5SDeY0rZ1Efvj3zAGAntouCJWrdptHGpR49UpMWaZPw
Rf0/pODzkJj1EdyVuLsFRfIcKX1pczeinPyqT2NvQE42WSbr4kt98Fj43yazDBETmHuctycbhcoQ
eJsQYIKC8XTN5Din5U7TW92BYl52pQT5AjMbvjkM7pIDc+bPLOwFAG7EwF2V62PCgSJiQKkqxFJR
SCboojVcvtJ0jnqsKu/wIf/Q2QUdKyLTl+3/hMyH6vULtq7L+sriThowbPIzJHY4tKFGKuGasYwz
uWtRrahwE9GHLIo/TkVjtNCnehEBDu32lLPBbsl4yKX7y9eMRZ9zqjQDIy9GNnLPxRCpegcjQ1Eh
MLjnOWux8bg5ATBpgyfWMyTmX/0P5VTYsp/OzuaGKYSkkVQx5n9PFFc371+40LNChT1ApS07Mcfp
9GCV+fIkxctPiQO4b7ze0JiEmIzhnDlrCgsq016sz1lKa5cBBY4WvaLhwTRuWOAbRxYpHWjO0KyG
2oqDZj/skyfB9nz6vEVuoagBkE5a7f6pmuE0+q3kFpcTNb4GQu/D1xgNOwCY1FCckOZW59ocGqas
BsGpS8uAWrwmSVKDUgMDMLgOs5J5ESgdErV5aO5zJhW5VzsmK5A+G5OKgx8hrd9O7umdT/EdNyfb
87xXccj8lHfGiHu7v/3aPDpcAsUeQv5iIq3e5jrmzLfWBVbMLMT79HVpsoCCsNwM9uXlxJqUhbpY
KeAF5KBXqLAcNGaWdK2PBlGf3PLlOgX6UkNJwhnTadqmBFdTGijEzx2FuXA1zTDhIDIm8BIxgA6M
LKD9hrr58lL0HZB5k0XU46/gG5w7R7ksbSxyIFsISdm3NlD8sGPj2ouDZ13DnMP1W10LidlgokMU
uyVVmqBSmn+QT3l96x5DCCapJoiwmFuK1oZyTKr25HljpBe1bixslXXFcGl6zE6/7VgXA0jDZgBs
O5cksDmDlfZHxY6etmthCaKj3Bya/eomFIrh8HBr6m3cAKzJq9VXNZioMD+brvIr9Kyzbc/wB1Z3
BhnlsmyMPHMDQAyW8Kb/u9uE9PTWIHz8hRh10EIzjUz+WWksMsPIIwgIUTMJf7QMrwfdg+qqvrux
dUf1eUPB5kYdqvH6YQ7mP1xtqr7KxcGJ97XLsOyzdJZGwLx0TChh8sr1fBmkt2luF3JdTwt1dcy/
Wp6rcPDZya0i9pGQlHZG0g/4Sn98rd11/s3TCFj6RUBDPTAxbThvSg/sCEyZyhN5UGLnr9VgbqBN
bFVY3bCaZp3ipP/b1tIHSSySYfM3Z8kJC7yBAQiEdb19NtXcKGtuU2+Q+QzFkF32LSwGNIokyGoW
AhWEqqWpEol7BNAm+gKYrX/EQUc7lTjMXyV3el/aT63v2zsAjQR0Dg0dFQph1MuG64dGBlfM5cq3
YXLi4koZSsA72W8qD/QraCvqHmAVwxgwt2PxZZE4qnmPqtfpuc3un9cP8Xk9r6qxdojztdmVqBG+
FlcyuDv1574/LOanKyNedaRYE4jdNay2RpfXdkNkp/nBYmMngZhPINFpnNHUTFulTA2CS6Mrrh+t
jtGlEclKfkOao4ckut1iWmxxtEmcxU0nVmf8kSu8M4HIIe5UrmSv+PV/DtxaBsAPKS45lktF7ntC
N+jbMbH3M/yVKVl71sH76zUkErhUjCkAZoCpjrA6ZbIktcrwXR8Y/EJAMfsEfhhL/HGpnj6/jnZU
z5U7G3dJUC5JrSzDGsb687cRHitTXX8VwhLwu7PNx/hw3Kn+ny5BeBJnfe+GW2VU2vkel6EVlX2W
8WxpX07eFqYYV9xVfw/AkyoTMv52Q4luQDiGZNA7LtJqNZtJjNKZtKjzfAicZ7pxSuo6dVwwJ2KL
yWhmS/x4aWTIO2mYsqtLBJdvd3L6SQ+swk/z2gXTlyLboenyl/EFJHQd+dRPwgw+c13sZY8r8+Vb
cdDoF3elCTbTz4lYLepawruG9EnJTX8D+2ODhakS5ZvCJZoyvUnEo7AK3m6WFT0I+6nqraZh81/p
z/TC3XZhwjevxx4/3/+Og1svjnhU/qwwPxsOOuex1lkqsKbGmX7hsjS7elBaU2YZTbVJ0IIPgU5U
/3xtDzizpZb9WwAVc1ij78iktAc0RINCzMn2uBW755NJaHx7ApxNGRhOy+F7V/ZHS1LZglPxhO1V
Emuva6OUriJyEhYoa3cJjgbkB5Tmj5nLt7Sss3+F0y4cCgZTkENtJEAOSTpoo6lHoOkAQ7J/m47J
g3QmqovYnROUvTBuwkccy0Ue4i+H0ltsVLisnOT76+8ocZak0EK54V3SPp/TG4btItpXT8Brvpre
kY1j3Rwo9hvsQ5ttKNOxy6cXld86nE7cbzqLyLSwxz0LnoDErGcLO83fsDD3AtC+59+ZgGKyipUC
KCtP9GnvrB17aMnIKdFg79yCT0VqKmQajTGCCEJmGKO9wi6BFpmniXQXapHeyiHVGAsd+LocMdiK
qLUWtk7OXCVw+mNq6TNwxst812UgN6ciSqUlneNqevcSy/pV0Vzpi8oXg6bAM3AHgY5C2lEJ+Cgb
uMwgZ9XTtNRs/1YLXbpndie/ihcB7F9ImHCfgrVaYNv2RFnHIQVSlLAumfh/rcjaKCbsK7b8W863
D8SDLby8+fU6HzmBoTR95pKOTP87Y6o3X4doH1b7PGMjgwqCT4glRFpuCiKLnQzEPLxKNxf1gdfB
oLQ8Gdh0WqWbd72CydM6BKP38zLzRvlSi48jGTFlV1PJDryT+wr+3vtOzkkR0g/l1P6bKmwdYTbf
hMImXwGt+LpR51v0iIvKkfDVJcLnZ3kemc0OAhl6UldWfndbVFWNt/xKZ6ZoFsjS68liqnxXXsiS
YLzW00AkkHg3JhS4JaNzm3jpq8hDBow11Pt+vSrsa1Fau+2QkeQWIQ/YkqtCB1IZ4pA7kcsAC/fI
G+ztfFTK5pYFpC8NsUBF2fk9UNT9y7QB5KfWkIQVcc/jXU/vWkBYSov54+/4eh4BIOjWJ21BRfBM
LYovBZpdzZz7GQCU4U/IPNcWSA9wMi1hZqRP034O4tdOsR9tVCVJHP1m5NlhA/qgfCddbkp0zev1
logvo7u3hjGht/jY1LKLFB8YmaVjDTb6f4G1xXtLOVSGuKYxFUsY4eXC/Z9JtkbcnuLUHg8dbdED
V0ju277Pd6ZNdFdqobGO79e91+Aej/ypNfLlHL8Gdrj8xV5OJJ6aS3nOAXUQueHvXwSCu5hvxBXz
b01ElYZ+LcsSpNFqT6S6hivc42UhRWmz8KmFw7OCX2aY5BkjdAaiwNPVRhPzWUYjuOzyRDFabJc4
ntSJ1uqEikJrTz+UHSVHGKWwC4FdwqoCF6WN+2ocHAsaF1FKrXY30hGxwuxXafgDu563idcF/SGM
dJzXEspWkon1MCBHYJkI0eK2HJ1wMH3f648vhBP6XDh15H0MVMUJF0avNDkzM9AP6WOhMfUHS7TP
Q3XyhRtrGdVEpMPrwzUdz2dnXKTZzcOrvbeNdmXXtdzsbE9MGSZBnalTd8grfG6/VJnJuRyUCNs2
4apnWfDPszfeRyZwQFed9JLJg3S6fftQAiB526uweTiMg77SMYZsFc+yayLzk4iejfLK6YNfe43g
BmDpoXU158yThDGLreCwclK7AJF+9n+TZF2PqgfiDvw4X5UknVhbJDw2tt46Da5dVsguKIYP9rNP
tuIlu8IilAUsl7n68mdwjLJNdl5+4X/Ha6SqJnshm2JFzp93fnyEU9tIw7yeKj1O43jkTXq7rfFx
7zjm5dxldYjAtsekiZCQWTn0cHhOPl+wh51PwP8Zk3y2/GyCjosBhzg52X+ZmgUtLZO1zgo+PBu8
rDkTCvV4DG8E55M8r7YLJA7Ndz77/jXDcyofrMSJ8I5fLKOmScjRqPfTmb4A7lQkaEPTAkzhj1md
Qgp5mykJFy/bOvEUJWmJPpKscPqsuudAFXZ6aksvsufkjMiwrbjkhrtzlOUGcY10AQ3MEVErbQrh
goglAL70p4mDy1MVXM9e/EvlPvE0o6Spjl+c9yzgqER6GrsYk5xCB+nV/81cYkqLGqwgnktiNdpm
PJhvjYsgmE2dylFK/bYyv6cOJGqXENLGfXy+6mxe92Uc/DlMm4LokFt0aOY+Y19uyEz8fSTlBzwW
fQDLf4Aa6A50e2eeBYnFbr0RVnGIRzXz+038PN2J7N7faWpJf2l2kEI3375h8i7wd31JAQa49m3R
9oswqoNU2c6uIbV3ffqC4QTYzlDL4NNRTz55hT/LuHoI1YSD6zd9kiaWvj2LiHy2KiDYhAwZEuCJ
Ge0G7LAhGAzkaUCAAOVUH7qOumTtMFGId+oDzrIENWU25bGCDBOewX6ziVZ8fWPs1av66RPzxghB
+znLcrhjotkx1n27qO2RO2Df1wqnMp6cFBsd0+fRN9mcWe8wZaerLf1Mk5ClWgHVyH2rZ4JLfrN0
eMq0mD9hFJmVX6RWKJAIv0rar3Q6tNfmQYJwHaZb18S8Ly4HsQVwq2kJ/fsLDkWq9m5OoY7/93lE
wZcB5rr8Fde1k+2ol8bgt01Vw5X6DCmkrMTsAX67xHjSrid3YsO+//aTgfYpvnjdhfZo1pN0E5hY
aGggZiLOeQ2R0o+qCfNxqHPwF3ZZVa5OcIHhSdlgeP37Zb3cnBE9ehaEuEL48nQjFgT9id3Nn2kj
VZjAvGGOplj79c241NVXULnbYpyN50Cg4cugJpO/u6XvKZ1QEO0kcnRuNT5APsD9lMdO5sDRNRGQ
zQih9fSNaSJ0kITjnYtyfqlziTSKahjHSL/89uMJtj8HmZMQoxXt+jHgW+4M8SWyejmr170933vd
PS7MbGSYjvOwJgaL/bBOnWD2MVNlXBJAsoAgWzWymfHBhmWiI2JnCFryoOBR6j0Jse7lc4664lJR
fM0EFw/yIvDWSMKsH8RQ0L4PDW51Ck6Z3uTUfAivGnaXm5u9WCBq+hKoF9pe5Dhpo2J1/90+O9xQ
9I+Yc569PPIaEgKJU9qi8frkLX+O8q2JKqTNQlMcmUOt29wHcavIxrbobRzHNMz7wedIA6FhVWFY
Zyy59oBrrxtbE/XamNBbC5r887UeOfgjbUmtR5k+hlB00oAX8PpaFYnfT/3pwfZJIviSi8H8tKrW
4RaP50/8qwbzqIpmhU3il3Bqr4lf3c7y90ryLiRu/bsF3bQEgH5odR+fM4pleSEBnIIIObnV7/br
SThWrol8jAver9C7Tj7qhvXIA6wDS2mQrh7CGiTlZIN1X7O3g59EQp3GepiADkgp18VEM8GJP1Ee
ajfWjC0cCH91Mr/2ht0P4148cPnYUNY3ViaPOSxqjRMoG7PJ+y2ZFm1uVqhfH+Qh3SLzS8ooVApG
7M5JzgGP19OqRn29y48sO1K3rrMJ1gJcRPyoZva3WCvsbe6ZxxRvyM7CYya8FOc5aYI1W3sDHLEz
lyuQJ49K3qzWUEEJ64hN7ueMLF6ZCi6eSJfDRaBoZZfHe4Xwad8lqumMY1gXBIjqNaFsnKwGeFGN
lmghn8fLCOEnHvTfYtBOplvydMQwZwQKmE6+5erHHcKQdOJRuK34AN6Dv13rNMQlc9J8uIzF6mxm
ZErGNQGXKTS6C3AywzkmxAmrtm9+3Bt2lnfXa1FzUJum3qudsbtt3WXFv8wWs7bOuLzCxO1FkSDf
/ZChNAp+aYlcoESxVDLfEf3xkLjjZZ170SeFD4TdM+gtpRWDk5ssWHLG/H5de3ghdnIp1XaLlPq3
bq8BPBi6TRhrZJ2Csdg0f9RadgOsEly31LZkA0mbG9i2cTtPTiF9OG1cyz2YQZvtS61XkEvNq9tb
tEx41RRVcQMHYxO8N1nceiXo5+VjMJ1/FPZpV/JL3IaztRgiLNZR9o5BBfwMhlVtMTCTUn+a71OW
/DouIKAtkDa3jhU+pEZvGvhnTBHTKDC7pmGKgwCLHor0Ww2kg1dqlUF06+caFpboVapVW/KzHtJx
Y/5Ef6ljueadBPGLFA2X1jJpLJwJ+9WCyNdzD6J0fHZg2UHLfuFJU7PMmAFh5fa5dwHHewGyEoV2
J9v5zUFCscfoec5zAz0dC9o12i6aTYD1wZI7a7jsfhjYAOI+VZiMUMvxZSDJHa9ejZrvotfyVDzA
1oz3op7BjEwx4F9e1e14So/QhzvZw2jZ0OWgMF2mPwBs5uwxNPWJXTNI7oprSDgtjNZnIsV6P0Zd
9T624svNHgGn1cihfyjanifIoR81OlHLQcPAMfkBTptQNPQwGfpW/nFDgBLuIOqKG7CWTMappEhr
JriamwG4dAoXrdBgRKsn9Sk2IyQnUvfRLgYRVRCaEkOcpT+W2PIqjs5KrD4F9q045GcHOZSVZVo4
YPVaul4PvgtFUZRzCg77FP/g0MSFBMRBbrEPTVwjuafvOiClsLQuR3rmwJyDisC6YCCDW8CraBcx
xlJkSLYdUJHyk0XG6lmF+E6s++U7pB7Fk3avB1IWPK0c7pHtb4R1yfU/5+9/nc5LGGFQSjSIX3NN
TIlKT+dFkdYAhR9ZHzYfW/AnuT4pmO8VUiNANsXRqvAnMQOSsmhkB1MJDMZ4VX6Mo5Adw3Z3Ev1E
+mTd5Z3Utup8ec830J6xy0wYvbO/Ll2jk13zEaCFIcz4JnM/DDkbqEe1KEhzMvOtYJOhirlKHAq1
cNbr7hkIVOnPfX731gCW8ktGIj54S+1/Y45AbBKNC8yf5TlIDsh3dnSiC481XQVz1RiYGUotflat
zug/QKSfCL7J5sELqz02QqD3F3oOw5vhROV3PDU60IBpIXcWb/qD6KBBdtvFlQbzDTCI48Bstbuf
92GUQe3cQx8YpbwQNIcoHRQnyupAV4oVOcSFZbOHaaoRqZp8D/ENfZe8EgllCGyiqY3si1OeH+OY
OVhytvQDcS/XrwjwDVE4c3WF3ZPkKQ2yYYfShIlQK+IAnhAsByH4HLIrP2lhjGnON3/BLcKiruBF
DCNscDaW5WneEV0u8MVDdhl7b2e0CezvD3p0lkYKLBynt7/Q85Xzd1AuvYrULT21bPwuq8YE4zL5
hh6FJ1nNe2RtnklxxUtRL+xmlujrk6puPXo0n2Izola+ZsKXjbAm1rKPzMpgTWILGW1HdNPhusJW
2a1HEsG2u2IkWGNRYs2leTl2xAxTfINli/2TwVG0rsDYj9CWtWK6Igv9OIgXq8kMOPrHw+24bklb
A9RFmm7aSFzJYlK7rJWI0wgzyhd3VT8IRUWjSj6gATXjp2I8ybx/FvX0/hFliwQ0DIEPQv5fNFKX
OyYdmdgaAEddlVDsdl5PsjVetNYgKdZEx8F7hdlV3Hp3deCw1IrGlXzN56fzJj7x3FzsNcT8yGxk
yA2FoV8x4NeCK5+3iZuccoIMGfjgKrNxa+VQG03qo0vX5vXquitST5FoJCBpfkXR6L5OlUaRazTt
fT2xi/HMUhdJC3uQUcJ8lAFsOxwzQ7zSPT9ymUDLZTucwljZ1hT40nsj94VpZn48l6bBjTYIGTC3
rLUDxGk0wkJ7lJeVrpfVJ+ii3pxC2LSMpew2gyWg3EX22FDr9oVYEJz9nhNrbgtNYAjGFUJP3MoD
1ZjkMwV/gyqSx/MW23RL4/8j5uoAp5I7P1P8CrkqMDXQHPldbvl3gm+qAZDjMTJp04tyV3IE6gF4
Uo4ccPl8sVHWVKhiC5qwy0uFgoPGsXxOtPQPK68zSnQb/eYPHINxQ4ueJkJNvPSD04L58SGqrr5C
horXL2dyLrUt2YHB+FatKGhs0yL321ZzgFjtp/pw2/La7n25f9r5LeRP/urVMjFJEf0hW8et006e
bkNuMNP61cyPTvPjF6Z6MVw7MbNCuKQ87SrA68Qzl8yqIRpGuYyvEWs/gvDUqQ6B7HcjB7Zw+4cT
LW0d0VL+UCmnnkMyonnjCW6IusiWLGx9r1S/DKYl0HyDBHF2VX6AoXMt+AZRzzgNA556nKa6JfC+
GuvffdQ2MhaUsYkKYqSbfI7vQ0mbnTGmGplL9xVJdBkxddbBZ/6nbnHWL8WHA8Br2bgDL7wjUUcw
IOtwP4Ag1Avkkqjlw37wRl4Wc6EB3PGRJ5hvVnaq2VQQv+buT0cWaErqsKKMZrT+bx3z4L3ZUDM+
/iw+RQBRvQMhB0bAqHbm8p7M8CkKZHoeRgxz6x5Qfnm6fdxb+X+jMc7p75o1ZYcof9ozjwc9HkRm
3QfjCOGUeOhegmfG2bjfeoJyTJS7xDEWfMk9SyODFKXJthwAByc6OBkDo3Ko0IHpEtRXxppR0wa/
MaD6QTtSpb/c456SBEOxbyFGqCRsVQCxllVqVakUfgyZw9UGO1Ek/8mjywFceFezm7YEmv3CjDTi
yi7m2yefUGKRNuSatlorW0HYkWeptMmmXGuVdLDRiKt07+cyRx/l8SA9GTcTv4tGFn9yhIdEi1kM
rzN/ZB9K7wLtfCd/IZCkAxqHIc6z2NT48plGhhrtENsW7X02uwUdKh1k/acwMJuKTNbtoD6f0dD3
G6kJ3cmC3u+Lt+ZOIlJu/QbzReJSBNHYlRk9oBlqvjoa9n2sBZYrMjnNnwdPyTEkNxxgzoz1SPvc
06MspOSiKA0nIfmXXmS7m9bY4GYqtXdvQ1HEx/P85dZtVM7jsxzXq/HCKPydsOttWkLWLQhUSTpg
1gkMHnfG4tZOk7NZC08TgJDygreREWeDmeShW9TpUglcbZ1q6ltxnWGe4EPvCFIxl1nV6Uozvxfp
viHxGH8EQir3GHaCQdbx5Xr79A7t5b6wirHdPw35U+LPQZ85uuabWCFVPJLTFlNgJsNEz0iR9L2O
di2naR/HGyHnzKydMTec+MNw75PtF5BYAi70K8hAiDd6Io21kbBBJOtUlAjyp6ZshGj0r7am3lJX
PXabRXjupcqOpeGyydkVF+jLggOMTUTfl3NKRXlqu8NtpMBi+WUKPDw3tcmbVaC50KD87Q6nQ33H
NgzA3EWBu5/1zwoBkaYau1xrq+dIbdLYj/jN4uLkvlpBgP1eqjPbTX7Il2Z0PSF7EaQ326jv/TWo
Si+2el+ywbNv0Rdn4hNdA6lJZAKXy29R4kYTMBvOvpgNmR4RVjZevpn5zGoaFK9Sns39vA5T+gDN
bnhEEuGUAdgejjeeZKsj39P7UEV6d1/R+RSYmuF+tFXVVJ3r04RIAKsv7Nd6FVbF820SPkbLZfrS
8SyNvjSoroJYKi3uQYsrXhvIvZYyjHZOmxtBT1ZH+SdMg8jmDbiaWL9aoXLoqbgCFve8L5y+Tg3j
4oEQOJo4WlR3EACAAD8bOtwupux1jlNhYPdQI5ZwF0sjLTTZ71j2dgO2dmPGKpvKDn+3A2bgwwAw
lx6oRw+jO1DPBPiD96TZRT6v70GAELZ02oVAuYygWg44SejSZtw9FFZ+M348+bIcphzyVbQR70Iq
D1PE81FeVs6S7hoqAXdEbFV39sdcH6vRf3lnn7gbCSorvM+oMekUCJFvyT+KYrVCvEIzm+UFG+3a
cff1i1InNsczysRVr0UfJHoxQDbq0wHZlB1mON9dJJed/f6spO7OG9f3V/wv+0SnkD73khc7f6lX
8DJXhyFnLbFtMO/F0hHjQ4/qJFPu4oRF8xTjsf6QKi1zTi6LV2pXZ4SW4exQMzjPn4jdMQQ3KHyS
SNH4LseElgC+8gebMaRlaXFAr9PmG6tiT9NbrfYdRQGtCNeQPpxKCYKkzYUmz0ICYpSwZkaJzVDJ
aOluhD+yEBjWYCYKlFTeVQNOHCmI2Ll9dS7YZ8CbBHJxFeLKuMJnswSI1cKcMbDD3bxW+yKAprWq
h4sPu7TZaXfYmSADscetgRHup+MVq80w/EpKJfOhCLkvjJMlU7MLGur+N9FIJ+oEBQXTEv259FHf
nXnmZXyo2GUVEUQ4V0R3xU52JHjjiCU5IIrfRK7srJWe1X1a3GiJ21FfB0FwrOWxIUs/PKmMxPWW
RcgpgC/C2wZShM81HyJlJ4ZIxV5mkkJ2yo67NnJ9RFbVYai2lD28ryicsmn2yR6JESAbwRpjqw2u
epF2k1RoRjvXQvQoLFh3VenuRxv6sb6n3+E385d5dCv1nhsTEqRctc3B+0dvr4GcApDLN9/756+d
1htDKxZkmBQNGrYoXcqudlQv7+oCJuBRFQa0wYak9FinoCsn3mvxS9UnHqn2Iwtdxq/X6P9dYYqf
CGtN2CqVmZzccW6egFrnGVpYAt6URxmmjzovfmeSwjJ/hLQaOeyxNigl9XC4pzAwJkDYrk/wUyst
CAggBwQYhLkGHgmp4DR3YBO+Uwv8QXA+hXciY2fEMntrmd+Mn7++aoUsROsc6rHxoWiBcIUduBwV
WIrUdu+gDgccgD9MXYDc6+w3c6RFeVS11wonzZyNLSA6QHR2RLgWISpd7U9rFoHcAAr1VxR0mqrG
X90ngXlXJzTFX5QnzcyZr6TRwUylo83I3UB8lLjvOKzc8aCrRixtpwltH7fgnAJN5+SuonmC1btb
sLW1kshnfkRur6qOJp2gLD75tZqTZht7vvb7NpbkCgDaPTyJny8NlRPRU2h4vVnHPPGhaNVgT4kt
ywEWQxLND/CXMGC+CDWxfd6COIluvx5fidxkwHySSPLFPmAM5z+7U9CdMbCphUHWSDZNV7BZ5W1k
kanQs1ko1rMiHAWRjJHZlZOqKyIJQDrFqkG8LK++JEdor+r9ApXRgXZfppfZVNp9BW9kP1NoJY/9
0uQqXT0uoBTu1qWsI6ORLqgrgncw4EPmNg10tU5rzznWCVdRGoZ4FXc3oD8sur4U5EY6mtn1XdCf
jp6L71OYztYhL6lzaIFW3JDoL7c5vyh9dWnHTpNE0xtTeofvcl8inK3NRHA+7R0KgS+ZOxRNGnpA
Dcq0ABfkCGyQ/SsFmyxhO0VVPfxmcMoGc5srj6Kk1g1SfI5m/Q9Tqfr3L3h9oCPrlKtgeftNsBNM
AmpVC0zzKGPchk0jYvT+Em/MwLbrMTZ5PX0JTLKHhfNxhy4Y5YTPpRwueiPtnydzYtOKFzC8Lvaz
asR0jzH0IxSVlcKcZ3EJmvzX0cjhcihtFfoU7B9uVbgszd9RlGSx1IHXYBuaNipx5y3OCEN+zJnX
UMwyTtUOpa+4MyJaVrLKIKq+HiiOCnBP4sWxj0t6uPevaOmZZCF4OnXGEgEDRQYFLuKzzy3nSXh/
fVSRQT6Tldd7GtiVMlSC5VXvMe48CTLHztRkRDYndWc7z1zIaVxE6tBQVLrTBhk7+N9LFoJNwfUp
Eqhsn+VDqWGN0BKSEArgXNivcGxG9+Y/x3bDB4MV5ayzxs/iRoOLs3xK1+ZHMhEbL1PDKFIqAlnS
hO1Bt2G78j4Xn/GfrWA9HuIbIoIa68RHjBTYbpvjeeafVpxqBJFpx+bgroYuxCWPYcKuRVnJB5fG
6iqUcs+ZmirWGMbHm8nj+lu17xDft7BlADSByuNIKmR4l3L4gz8mBX0kt67PZdK2sJP3nMVx0aE7
Haiu39d6XVr9+2lkFMNg8mX8bu5369YZLL5ok0Ks4dAmuh16ocFMFuXckcY/XKmpIYLedI8FSoZy
KNUQgiCtMi/mhMESu0rRvxGhliTUkeFzbUyeyPTZaFJ7Ge8p/CJF1vHYFSQCV9GOyiDMShHTMuBl
GY439Rp3I9yyrXie9/9kkz3NUH9ryMGvllOxGAHLuER3T7RJwSMi8KUeqpmOOLaGL5jnnTw8XRhA
lAoIms85Gej/K8mJ24g4TkhWtPB1ja8EThgYrcJqmd0h6RXsNClrkmk13kzalNYhqU+t3UuXMGH4
FTe9EA2EcGgg82IHe3Omvza+XYND/eyC7Uw7C9/zMCLzT/Cvn+TRoSJa0mZRkbitlFiZEmLP1YXY
YkXypMoOjny2kgIvqbpCMMsYX+VjFJCbXfpcdHi/W4c/1Dck/2au0sLDGUwx5QSiLk4+IIHDMW54
chWaSiTeDIqT0/RasMO6RfdDwRxW1zxsAewejFaNR9JcbckUlI4ti9I0dsGFBYdwkKNfDWmg1MBh
uMklMmbrOGIFpBCslau/mXBd9L9SMOBJ4yooVcqVjCFhMX/YhqxRwueYuoYQ4ywr1/F5BtIuiMpH
mibAt2VtkivS0vkdtkzem3B9UQUeHmAvCuFtYt5TLyLlEnocHNtHVO5sXYCnvrf/el/3FAyBqrPC
ExBX3Smr4hI9iSCjfpftDI/1MeR4FOHVJ80pPmOPXjdZsn/fLUvrCitwa88bTSaRcJAL8YHSJQvy
6RTAU2ymThM65l0NFYWGZy3/d8O48Bx6qI973Pz03DvI7uzsoM2/Ovwxb5HJcvudqgaRCIKagGIV
sAGvSmv1O2Y/PzZX5VVJAVKAl0yy4GkmfKUs0BBmPG5Z4t5yzcbhUYaOrW3ncev1WITgpmbtae2f
7JHasXBr8vkIqyi8dAXSW3DsCkDH7bSqDMUX+ZFnaJtM0a+vtqvnk2a+l06j9YVmHJzakwHrDE3H
f4tT0IYytXH9Bq5AzhsWd7njNlCFIfluAh64dGdoC06mFKUFv9mfbQswWb6Bi7EULjm6niJJrmOT
LOr0FSJ0NnIutlbpxsuKYZvkFMMz0ycMUQJpyS3gfLneUHuRJvhBu+V/lli+qrusFcw48zcftXDX
xjaZlXdd0YKSMTwUf/Pe09+SVLBYw31vmN9XYE54f66wBaV+VJArbui3X5+QzhHfGJbw3a7iNf1c
IIb0w0BiZr9ke3b6D0ruhiNLutPSjkt50m8pXkXjKHIFVZK0eA2PWK3sN85oHG04neZOmv73sE4S
5Xru+EDtqsfL8/oUmWMFrLa2ddliHASGAYTZztiGAH7Px2jas8bQf9QzeejoElQjHX4oNE0AQERy
hlI4tkMHcRPquSfNOnNtMltv47zTBzp63tLvqvkpqFRaVWkRqaexUW0P8pddNp8eSBAGO6/Ttvb6
qVki0JFk1ZaWZI2nJSeBzenw+civ+iHO8Y/ROteNMfgY9mtlB3CAHCpgedF0ZmqT5XZb/bgKYaOg
tK+fGJ9TepxT6DZ3PN9ZOc8Kp2DnIK9g8oi3zVYoxaE0FpeVQRm0h/fOMj21hGURo9kATmjMCBGP
3JSXRRw/XnKQ1RUSZpBJgvOdgBeIWOQJocXK52oVssHjZDz3bjJ6KVaeuU6zVxmvZQgMpyQ6+FFo
WIMnEjq5DBNZTiCFJq5m0r6h5dDGglfY4F/0uln450YHEulCEhj147yquxBS2aYlqZ8LOFMH5rEv
rbuMaB5X0X3itM7g+pmuIc1BRCj2lcMpCtVdoOCGHW50tEFNoWQkNLB4xbyZY+eIgtfLv+w7PqI6
PsBbthL6ez2N+wACuY+TCQgzUdVeHvp562zN7uz0dnIv3BNR5gUOZxJd6cwLu3aapsVjLZSPzyav
qkr+gkWyZl0a/oCQ6JyOEearySj6jruocSFT965WxuatqFhc3gEZfJzkGid3W4ujqhkIEDaeYS+O
cBF/bxbLr8ybIXhXNpXuh5k0bPeMDf1t+vRjKH4F1OEHOb+uz5uQvz0sorCkfskivKVDSnMI1oNP
n/zuN1RNjl94FSRUgrXr3q2Is7gO9R1m4UIyYmpTdKsG9Q4n/3dTacfdGniNIADzDsgGSM4opTJe
MwPFQbhTneCt3eZFF+rwPPXDuQ6aRvId/o7NuTbU+qBjx13SB0+KQKlSP8GBdU13+4LXV4XykLzD
mutUhranmYOMIapWYXR10PFubOP2pND6Z/CJd7JBzLFgmHVZE/A+MCqr0YhxtNYQQDhEDpCS2ujQ
oPurQDezDFgukoxr8MEuoj2otTUKIccC+XnxICcfPqaTzJiKwYOgBJmlaSpoiFAGQG1klFAsB+/B
gr/QaQmkh8BB/6cY+e3oIthW8TIAzc77WaLHUkGnESjnCepXYobwz3YLWmBuaQKwu0xqHHLO/nnb
Z0T0/gTlsMNfJ+kDZx9rrWVdwe+H8HE/7h1cFNt/x4mOL/mXTwBLmpLgx09/zKb+fENk75wN0Da6
MkOXnsDc8yqpxTHDOEl56cWj7HqncUXEpWK9I9MBh/cXHsRVZRTR78XZCnpjaYHg7HK7+2OQCJCK
FeagYgFKg85u6n/4chkwNrW8nKv2Y/ml5tVH4u28e2fhL8DSag6F5j0T7IyX4P1FJkIIRM1JrRnP
F4ftEQp9GJgKHixx4EkGAhghzgODbZIpar1jZpbvXm9KOyr/biQikymp2ErlqzzfQ2a+skgqfhTK
rI3KLOP+S/obCNXGF0AmUyad42YLEpPF2YBzNl2iHjIZmC5nh3xKBaHBQkBDmAY6JlAnpFK/nIY3
9KJrSfaP/1tT/TaPJ7r+Pk8UApX0jUndbXUs4WRkOeDglN0BjEFlOpLTrqT+hYSJKD6YD+OcfLi5
Iw8OQKgnnWS/Foak1ME/qXirPyTvqxNFvedXXheDXrcIziMqhlG7o7+GVnXt40WmNIVbE+NaHKJE
358qIejFiBAmBDOJV07uce0VTt0rUrrumehGWEpv7jnibVgEl6YoQ0YDx0bbH/aYffl0Bid6zOFU
frnVCAkH8ZdNtw8+/YleHWzi5RoEFMOr13GvUczvcAiy16fvOtSHAjCDab/jqgGqjMOb+7Ia8F8d
onPC5M+oJUcY8aQcxMaiOPAmkjpyFX/m7fpIhszn9g/Goga06CGy/4UZqyCo2WpmFVI6BspPXNq/
dj3IGmIQ8hYG/YFV1rGzPggf7LyzzpFmquo/4ZEDQ+5k4Tq8OCjkvsW35fjVFbTIND0L1eVMVyGF
v4mvGQWaS9M/QYUM7mlvGP/0e4rjie0Pv8gdEis2l5K/UjwPV2zUdxgGsmoC5OrwV5cPVzAs7Ina
E+EEXgK9Vxt9LkZ8Khw4adJ81t3dPjnHNOFC3PaZF4FkKhBNL6uRGP/OVxabtRjjEboRBK3u2sAy
oyhHE+AHiPJtBF5gGf7pv5LkF+vh6Kz0ITOZUWpOYdgYiDzP/0vob8NbgD7rBFqJqEGcrDRB+brb
rLu7Z94EwQOd69Fh8Bn/DMrOfUQXK8HNveeYvLvlQ0GFoLezOG5dv+X70L8EwuesnFuJsVDm+VP5
07GCFR/BK+pTRd4UNmSVa7pAoXncarWP5e0lgOF7ZJl2ygle7FTGjNzNSljg+OuAFDH20zXle4E2
8oCkjcgp+iaFmR5yy/XeRe91y1U5u1tXpYZy6S1ZOZsTaUM2JoWm7dAoc3Vugmxx2CRpJOOr3fgz
ReP98x3qIxwcefoPVMaQIALew/vTtc3y4j3dT1lLhinqoNf3V5Fa118vC3hhQBGTGbj5xlZylldS
SVJgVhSUbzqcqJXfa4GQf8a/LpPCfX+6feU+92Ko51II1Rvd6Dho/7Uv68xvofTSAySoKCAaiMCX
enzRSG/nGFW/LcVIGbRfec6EVqF0VupReKROIvMYc/6+H7elSdZP6wUEEsxxLv78phqUCKgYY2gk
C87qwlV0AC0yIuipj4guIYwbuJTmLrtOtVFLl9rc8k6Ml0r1o+FoVYC0tj9O44LoqWJWqVuoZ1El
LSP5bDdGOXWHgTCNKSaaGxaKYNjUiQc8Xhpt3tg+3EBH9DXxPhY9eswX3LMPxUYBwyjeG5w0/PfO
YkptTybB+CXjlklMexuM9OT1ZPI0Orpxo9ODtUoyeHimpXrsDK/X2e+623HIV3Jsj5X6fzw7vDML
34G5x6xO2FKeoPyAcTDjB1Hp6LATepJ0q0lsShCoaPX3jVbKGfAjrHtpQw2pWnRv0wTZuVTzUFQd
LeLPGNQYpqAbENLqUNqjtp3Tp2bfAeUR1zd7jAVjvG9GYTgq9FQQYnU8azDtS0IxjmrliF3PIHUV
uO8LqkUOSolG+NVUR60idoZNh7STpZ3Ys2d8lIwIhzuuMlN8J2p+ZJxHJz5OOcsNwXwoS9X35HIC
rQYhj1s9SZU7CFJWFgjM7bJn5ncxEbH0BC3KXSCcr7Z1QJ8j22bKXUYkPsjzlmUZOlwHhV0Zvjo8
M5XMlwgG8bbRpfI6hWBn1zT60335e2e6Kwy5M6olWe/GpKiRqotxTvdTVD5P0UZuKcgMAstP2cPH
7BWPaZBKyU/IK8naDkhUapcsVy2wwv8xDOjHkGl6zR79LFmyxu3pZugenpUAslJ/R+PpwH6rJhoq
aplgbOxCaq9p5pLluU31gfGZmnBrcaPPozXwT+7A6GMnhoj0/KzAr6zyr/Vbi88f4+FMoBwUkJK3
JDXm1G38hyJFpKksoml+as23SpugQYkaN5Ny1Wzb9A8W3v3ooPxQZk8xMDQ0M8r1152odaQ9csNf
V/u9ebassX/9JBUj6N9nxd9119zOBhwpQAi1aWxVccGqj6baTIiMYt8xMos3tu8YNUvJD/osh2yq
RbsOz4ynku8xB2z+seAlDDGJ6NaUQeL/ABJ7rVojbPKEQeTZv1tMIL779hATSszD3aNPyAoR15TO
zVtEchkIrIaD/qoLy1s6Cw+xUinELXmTHjMRvE0cKEz/qd2HZtucERpCihnK6FOrB4YAzJ13l1tq
SMEbXtw5MJa2FLJ3KEcffzyIb0ndCxrgjz7HvQ1N5qvCHmZj/z/MuXKYqwesnrS0EnwuBw+1PuvD
65OXc0j/6Z9kGR4evpGmvi3NSd+HfXQBUWZgjaiByzsk42DxDuFTJrkq+o5P5U0FyQHqSdwGwg9e
uMKuhqDPNRXM1dHRzrpB1gyQe3Fvs223YQtdDpfUsciV6mkIKJWB6ENiEBVRHAYo8Y+7bmAqorqM
OLLK6+SO8j27etgyFABc90557yAB68wnntF54yyM2jAVuYsTptFzZxtbFX3wH/xgNHga1YWxMlz+
mpllGuIIu/WSYFcZHDpIjPwU/bmN7gvtBehfwFUUzsbm5ceraLy5XqnsmHd8y/KcSZ5aS0pNDTOw
ycBBIif38bzAm+wMbcDsQTCgRLTev8a8lWEeFSyQRNBqaF6UWB8+nHkb/Qhdls+O4ffIsEolncw2
pyex+Rs6VmyBeVUXpRDGZrBUU8J3qwlM1yuFg5CsDQpI8kOpDynYjEvulo6ftuERVO3QDqFEOBhk
GWMamHH/HYUCGkKzRVTVumWtwR2dtGIDXm1Xw/woaCN2xVe0wkZ9sZTCE9HcmxqQAe9jzzFLO6z6
C84EKj2kCmP4oqqwYTX6uu+bMeMS6dw5EDlvS5q5mMEzq+fMIhDy6UEvFqPBCsT5UHCEDysAJJS9
JpQhM0mnAISTN4NyfLo2Pb2zdWeyqHArTD186ZDbpoZJaaBgqzM6shGRESd4UDVxP5JySMPtOvrV
XnyUc9JCe2d1dh0u9jL+MoSCcd1FQQwflbUlm6zva46TaW8rPPCar+tk3DCHYySLhPSai34DWats
52X8lNCkUjWhpj4q5OQ7xw9hr/7ZKEVjMVn7nwLchBC1SC/P5EJeZFvEhOu69pNgxozcJVV1Z81l
9Hv/K2GmjuwFxiUCnZu7p/bejWRKkkMA2Py6YoOLFBelInucjfoPUrtycPh72D27PLhxk86hHCTU
YzVYX3+FdiJn++rvEXzndIsjNGP30mBYw8CYXm/hpeeK6LLvnibv5sEYESour+uN5hKZW5GmTABd
nucT4etMxP6mohcInklc0AiK7w2qf8ayAVXSXOZM4Yg35U74wE6i1CuVwMefymnpRx7J4PsJBNzT
IOaHvmW6M39Wse0AxRWGokMnZ6lVzuBBQ3eOlfC63wnuFbpVf2nZlDIHDfURi0Gg2aep1Z2BWIH8
jTA4MMz83Zr0kkXbVkWyuqkctonIeHIC3QBZhMT/b2p49PjxM45P/TUHB59i/XcbXHdQKkOBwg+S
PsX9RRxjKQD7niJiBOBakVP1Av0Wm+roSgYV364Rloul5jqSc8UPZ59jox5TQf/h1T4h6UWzgKX2
vtdMzrgzj+kwtEZ+JLr1HOGDDhZ5sourjjNPELLg+aNWaV90IxCgxe+EALCJH6c6fcdPc09Jlcik
Afu4LcMhTwOSjujVJfJIRJtgosSsPdHrjlJUPzZK95SwNw7A2CmqhiGzZuSMQIJzb19gRnNJkeI/
s7twB1Djy8Sxilw3iFHywSXWXLebNfyM7E3h/Cuagz+YW5ab24iig2+B00wtpPP48c9WVQwoPKXP
+CZu5QhRHFhrSRXeUhznErp/vdjMVBta9/IqLbcgJwgHLXjeWIR8OD7UJpoTuMMYkZHj1ozoIUBP
iWAemB3jsKcHLa5xIL14J3DtT9prxva9wD85NVlZzHLBkt7U5eqBg4qvUeHyvDhp2OO8uBQPl3K5
yKw+cl+bK4lsV9b78PoNbV4F/5H9+iAPDthVk9PR1mXTwQ2bc1a+qWWj55AeQu6o8Qo6J1sr9KWw
Mv7eZPTPKeLIfEd+ha+FkyUBlrTRFUt7KByUOGlXBfjb2cjyC80Dn4UMVJsPhOFxg6p0XYIR3KVN
SdteadT0PgnZ2PxiYU3zlMS0RJq8eGUXG0NrW59OifRIiQRF694ZGwnyk99WQ9Fd794Mz0ZNqe3v
0jOmGXLiPbs58w0cQ55eUW31SUzkd1/D4jdgJB0DtOmZE2yy5tD764dbVKQlC2ks7abURp4L5Z9W
H8RXmHOEAtsdT8TR+EBhtZME1UcrjzP0oQT+9AOr5I9W6VNu5o19nsNuaDzb6z/iwFcgxRjjYs8V
TD+S2X4T8ABflNbZtFPJtspVy9qEvReQgTnxCHXIWAiGOwwQfSyRdbZ3YLUU3ROpBM4RLfW3y9m4
k+LhOdJPnWr104Ui2QaSccmHbZH8C5eD/Q3CD9C6s1jk688GQslvv2qZPt3UjMdz9/BizTbHwsF+
0avbnqcufVWSd1zk/VGajEYCA/7jjHAWL/BAAVLUNkC3M5vUqEFJX1RocUuQ72wP9uG+bSAdzROm
5vsoQp856r9ul6T3Pj030suUALGCqwEQpnzf0gsKlohZ2mrQHZuyZw/JkLk/BgCMKciQet0OStid
UrNwEmZA9u3rEOxdpUcNGcK81l8RZ498iqMqKNCeIUDaMSk/xm3i3JEU1MytRU4j6gUgVH1jcYzK
8nWA4jmY4IaqAsFouRCDFkCbtnD9b+arSCc1HS2xQS1p1Chr9ya3FWvuH7m6kHnYV2/utZZNHqKR
E83RHQMrf2XLoVZhvVWfDCmdxpzWOj+aT3CqpW50Y0zlxR1M4Ul7dZ0IeFzjuFxMBrbEb76au/ji
/YfOwT1qnLVOTIcDrIWibbqH6qbIHsd/KyGiDJ5bEr0HxR+fZrh/pFtVLPgzfx21uZIbRtmFw9tb
R9eSosvTIlY+z9rF6pa7WRqzODTypl2jY4yMCyft3ETWVtDHf/Mho6/WY9yJdnewJpxH06CWTrb9
2jtPN8qSeiQolkKGINpaCscy6yXOb8wkbL77gfnjtLlSe39R+Gq6ZPf5uaLetq2kKHVVL1P2MXor
0INDm7WNKC4mb9TcUCcoYoZHFmzplcWQ9AqTm0Vp8sUyVbvisUMkyLmvM3Hs8Inzn49c8Z3CQaFS
fAmrUZhxpwM23wh2j0FGhk2VLpNWMZePMXHKTFw9Ab3b+8bZFd7ykuCjXC5drzpmmnT9jsikbzQ7
w9T+d5a0zKlDqfbA4Ebi4Vt50zvrkYaxXNOfoue6z0ARXS+4+F1MP+AI/qMCrEd6Q+9FbptdZAtT
MdSWbEb/MeOMGcTCXYdutlRpWoUSGh2UKKv00nzTqmKN3fXUL4F6ZJewmAEQlYK3KBno5oTwkEHX
buyTdHuPSQeNeHHUhFU7t56q1F3TZ/cZul+kx+SIX7JzBuo6PoZw5/9to/4v+rS5bZrBWqkm8IV9
73cZAI+CRT9KB0SFtTWA1RTO1sV7Y5OiGEC6GCGLRa8pzz3gmIx1bDi5cI2UEqctIRKsNDuCVToZ
/7EhzvWR7VEuzvtFQCMOrVEWFn/3h8TimoNYw1lQ2MZKsvrBUJqfJqpBuVHSwBwdq8Skbphqpd14
utaOycpbthXO0H2AnoN5u440ojAsv9P5jf+XIEQrHvSNECBgjp+1L+oWc4qdLAqJmGIgrk5CxWIB
9mlbPdXTd191OBXkEyt+N2YDfJLnQdGZ3tHEMqgA3fadTI6ol5XC1GI3DdwIOzMBjmCbO0ndCVL5
bkaLkwxAoF7oy293sCbYDYu4Gu1R3up2HpEVz+PEQp/m4bKXrsmkbMKQffaFXEpe3PEdHvzXhu+l
Hmg2L47+eDMgxIrfdiWRhMCYC8ALQppp8T4DRUi8Pay1vdXmX+MQpeFK5cplIz8h3Pmf1wwCdvLD
g37E2mWUu+ZzJIIebKiukf68QlHM/fdSroJq4Jxyl8BBwdQM1wqdy10S/KF5EDWeSB19e2i/liza
OaZU2TOcrxmGnDnx+f8SpOjpTfygLrf2iMeMarzgAr7mWqz7v4J5C4IGA2NjFd0s8Wm652ngg79Q
+jgE8GUp1WzKVLtPqjCG+qlSuh8thmC1SOSRcJiA3fbOP3Oz6jYDLOu0OVz5XdY/LgpsN9FzMcZ6
4+LmzdYPIWl4kTqiE3eJ+1riSBVQpqCM2K8r+Drd5OjPff77QCCMiYDOn0qkW2okUxu3JtGJJGJZ
63ajis64NCi8gJRwa3HmHbvIP06HEt4okrM2TW1XVUMc9PHroYuGwE//sG1O65ro8sZNwXexhLmB
KnCtDthuKKQ+KEMVcafinAiqxQjB5U4MXlcZpgrQpSDAk9PBXTR2hp1jOvH5+/8eZ2YZUiozN/Ds
RtFRhLBvzGCORIxDXODmlU+blPo/2q5l/ASHSrxsFVnujbOtUt0rWUOrnGbZoG/3DaTT5znvhMIv
sKlSdRE/kwZKgYnbf3YYQSacZ3Vx+U/hUVNCkfSkV4VO+wVXUA8uRuWdiX4oIZRq/0Bv0dFkccym
UcjzsIRBDOCrXTR7CJg8ytquQWIP5ZOyuVUd+9RGThc++LoQ3WwJudzFJVbNQT046aHnHdw1vZkl
c0h+TqbIonar9u2uT7x4hrbytnOYauTOlv4YsZYTuHX/T1SBsy6mM192w3qNulSKXA2QI2mxMiCd
YowYctvdcVxsNXPwNUA7vUH3zO0JfIuBB6HCY3GDHofZXUrorZAOStaZA//RidKrLczxQFK/VV1T
WizmOjus0nkwJj/D+R/2Mv7ZEh45J5iXYPlV1XYQTWQkVKT8YXIqZ+f30bBqeTaqsSVIWUHLBZjE
yRlaVaZ923Z9vDv76RruHogioDGSCy4Gmjv2oolQhiGxqlpn7FYDEIuafHNzRwCG+LTssAxG/qQq
MSgipN+7jWjNdSfa04G6QpLcFWcyfAAnyEebHX39C8FrQCcVsaJcDgqqYgu7+Jsf7UAk29sfly7W
sI8VWqlYUCU/oGluNgjfcKdbIbWGTncudZtOblG6IypdU5R0pfKXDQC0ckCryveYs5FkFFlZLT2x
rxWVYEsWSiq+NBGZPvb+L0mXOwmYplo2FwT7JU3dh/hu0Koig05pY65vadbDDa48lPPfPgtrTSa+
m1kAlR8EKlMt4REpM8RNX7EvQPEXsKSFhqmdmsheTcyrwYALYjd6heBWj4FMrVChE6AMDyPUzdyA
sE3ewSepsbJNrMeCmmEdKlblKYZH+gvq0Ing3FqAPjdBbrw0FIfcZqu3dza8Q0LScXNua7B9a6g+
z24hY+dkRWhJSlCo/fMomFDZSC0xVtUc2EHtzVgiqGb3Llvol5j3ByXYhxxrVfmC1EHFV0pxpSnY
6ZuIO4mkM3cH+pzbym5YZLeFAo/f3JW/vmBs47ILhGyxzNDfNhYCOpSCc84anqkvsUnTXET+5yol
rRpZ16vSmJIZAoNNgzBEyl50Z9vV5fRDQSmGusvGar0RRx9C89A/FxW5zzlgaEaXm17p+wTKEptE
LgIdvm5pRAd9bRZHVt84C2hXI7we7tKApuAAshfPq8hFmus8rE+eXsh6ATAgNBO4bRfB2Qtu3zib
ZjLhP7ffEJz2f3I8yCbUwuWb/w4PgBm51eO/2Y9CEsOGEbpNusEnSHUhc+Zfl5hWAvzRT8wLLDHf
5mijAQIYC3kHhyWXm6G6ZA/6iVY3+bS9gSAcSNUpSNGAGhaKaM9/MmyZI2gy+skiqFErEu4vvBO2
xxWQejerq+Sjmx1q+zVlDgZJW5sAv+snmiPzb6jII36+8pc2C7OkwMM8QrQpMun0tulrsiifuUH6
lwjD9/zZ7T3Gc9XrgaD+nvv052tmqzw5/JvzjJR7GNxdLTwShYRBrWWI+9FjqW3HzQqH0S6K9ljd
CGfgCwcaY5w2eUtiJhkpqvGIC204yap2epjJ28/IRo0oORdBeuWfPKemMgwfeVrBhtZwy/8bGo7T
yIax5gBhAehoocdk686BovoiA9nmf9fUufL51C9Ho1elXROHgMrq86ZymGmBxO1d38IyK8afRm3F
GvyIxZVAHWNl0H56ZY+3uuhZ0JddThCCOkPiaayW8JfX1H0ngiKryG5a3vo8UDOt8RmdJoBIg3DZ
Ap2y+L39HTXcb0hi6YjDxmj5Oj6NJqBQjZnG2sv777IIS6DHMucynfVDE0JwGULv6C8Vu5J30DIi
OnguoTCbJP068R9G2xg2kMrROVLBKhwp/tbQ3++jn8RRoBKgIndrBdswghMy7xZsEVmtaTbPjVdR
ir2MAtIp0tFUgzgwRjj3gHlDP4Df+VLYdCWOZh/Gph+eHe0HNIWKugHhYKAv/StfpMEjtY4xZTzF
I86sw8fJiay2y92eILW8sIDBH9sBGriyWKK6JrPpbVNLUzmILkttecVW3pdmmdwMlJY+ivJT8KjU
CS940VniRdw86taQNtkC2VkOJVdOGJ2tU5H/lyZtQRlUADxUHGMJ35/EQe7gWigVuifxD5/fAA9d
sczU6a2/VXhM8hdjaHdm+zw7bMr8/beYqVxw/CTHWACXIUfPfaPkNWreQtUXee/eZqMUsm7z+ZZD
QcbZYu7uDdX220J/11Vn4Geis8wMfXDqget4WkhWWNOO/bgub/x4qL0wyO8MQTUrlpWMKdMZM2Xt
xPSR/sBOP9f2EYwMDHmobl2oVYtiSgCNwkF1aVkqrkcPlf8Z4VPuVl+IvL9O6rVA197U7wj5FlTv
FK9F0/75mPr/h2TyJMeh8WU27YiEY8AIBVJ/tlJx47btVMmA0vQxZ/7Olz1knPdYX4mu3SSNba74
6kaBKg9ZcSquVInv8UUHRLN/ZuzkFCMrYQiI+uC0MWWq0TV4AmVOqTR4QUi79XXAdYwrcjHVF+tj
g85UXMkhmFjryxf6ExW8g7L1K2WMqxq4J6wB2UokLPZTs4zLbZFL0pwja17voEWxrjYleFQ01As/
h9ny/gMFdOR3p5wxaTtrXEFP70OUZUMMgDSSI8akkbLEtEki8WEnACV+8Y7iyIfggqtjtlamiI1e
IPKfVeeAGbLTGXjKHlAsDGIebMSyNDuqgBoEsI4rr9D7yZU4Z7rJNfJrMXPoskO2Wl47W0G04Qq6
MTKesCRZ5d9Tb+CGZpmmM3JjDUQ6dRsmpCPcmyl++gbyB2zyopURJ/4Yz0hYCdOvwaBErDvU3YMV
9cjT5l7j74RGPC3+HPALksoELRCXLCBfzWxYGfOowz0usqphXDRixRNvsf8qwzumdOrEGhuUDE2C
wEC1/tM4QkClGhXhodPAINI9/X9DLPXenDWL0TV4aRRjHBtnWidY5ady+pMn17cY5YdwTZpQxnsF
0XZar3tgfAS1/FpBpauRS1Aw5FRLJFgTHO1w3X0FHRXkJPOMgAjl15+Y9YfKTFaDvN24G8yYQYu1
Nyifz8wpah0CKwhl6hdsOmQZBodKxV92hwrgLQOEO/ZHmG4e2BMeRRkuNuVzhsEb3UurjP4KhLQ0
MzNr553KiQUH/TnVOKxdc29jLXHWhvKHl39LaUuEyT1bMX61bOTUbIIQXC3PTitvk5K45lQ0DCFo
uB9SVdmz7UgtJICpQa/oLoGoH+C+IzBVAwAv+IMHhYr8/5d4r77y0zr6Qc49h96I64a9WTLGmJCJ
jnCpNnKIAWb4Lgyp8K8L3LrHxfTwEGx0zTfIXkggOP2mFKuAxLdG4FY2DxPSXA4XzyDF77NX7Wno
P2imlXGwHay5TwBPMqqO43vZY3TIFVtIe0KrI1guYnY9sYdMBIgTVS7bDiGq19hER/EWXpsPZWdQ
5mroxavJJ1sqN7wPUABckt+Y9uZAHDUdw4EvX8fiL6hwAZAfCBTQp/edqOIJZ7xu2qmcv/g9wwg5
8b+P8cLVHocADcgUlLGDfn8aA4+uehPHVafMg0sajBPkVcholBxs7Gcyc0x2UU76wyTRJP24owej
aP3qW4XAbrHVIDVfIHrSFYGkz3FNeMs35hie4bQnYmtjmxSQ+2qoIIcEtitKvyJePYfU3W5+1x5Y
aDbE2CHuMAsLYzbVGRmLC2FIbd2oG5NTVLxrSpYfvaZQCNqusMQpS8oIEnSJtjKwJ50G26wGoPOm
EyusX/IYeQLMq+ftha224PtVzrTJT8pNFET0chTw4QEPSqkZQpSowQj2jmlJwRHn3VheA8cTA5Ti
3hjbc2kfLy1rsXRCiWwxRW8sKIlozKpQegdKF+1c3BjUSSg/YiKtLvuvfVOUv2WrCSkQ3mzfrEfW
//15ssNQPWLGCOpTDRSFFpojUVAKNhGI4FlTedt3omGriFuwO9C90RLovoS7YvHapsaKjX02aVqP
XueIq5fWmnsRJZ1h64n348n9ClVTVOmDhqzRtcIbU0c9DJq8hNKgY1ukEpMtElIlfnLjORBQWor8
pLLY/zqT5a2RIQ0zU3ZWQ3kcr4lP7V9djs5e+bCFS/ACBL2CrUNKEgrPe3VW3k54j+Bd+BLEEl0J
TQ/CmNGDRI9tBWC5bgfUlNnGtd8k6kmazkJVBrcMCnUKn3LqdvXr8tCggj8brW0YLXdDtZBvReJZ
fRbZTYgcNaDin96ZK7gUuDucL4W0p9EOkClIWVrsLOJQiak/O8oUs4y0M6Gq1sEcxdebQrhh9w2j
SvObJ6EXMi64lO9FqWeYhDKQelXoDPRqCZVyaneQcBjeZ9eAiWhyQLrD1ObbzDbqhtOs6y9ACWQU
DOxHSs9U8LLaBZdwQwU5A9XcKVi7U/gq+w+CT9k1UAm9E17aK8eI5dD2tINKcCdbGZ7hO2RtZciY
JKg5XpWORA0KR2hW1kxR2moFVivZIHfCYFjljncR8C0ByZ2ftWcvwFhDyKiUuBfo7sxwEJfhkygn
K76U+jv/VLHq7P+7+SIYpHyWSbGSc9eEkU0rLLieFlB+5as8e4Q4erRkjWlUrsGqic+KcmgLWrX0
sqVUETc4x0sH7Bnn98ckUrrUSku00zRPO1oGf8jww3PiS++KwG0ggy6Hzao+ME3DC/N77HLsiwiR
ziDv8JrSR4AvvlBEYTKXJP6IzjDMK5gaIRazDLvHT+n0AMa3piDTKQxGRBaOoGHBACICmZmXRqDQ
i00xD5BtxTmFzU8EKCKpVGQiOhXP1Ob5MP+xAgNr9jAKxVKv0n6rKamVbbFS1ghC8IJKjxtxW8Tm
hi6HILKaF6ucKRttTNrkmQfg64nCDCb2EknWmwU/HHpwiHyVdOXhPp3NCOhn2MJyOrbQz+la3C6t
9Vs5D58y3RjN4J6Asd9Gbe3EujZGGuyWyckBqApF/iDI/TaY1jlqZHDSPGYhB65kBrj6rJsetqBf
3EMkVFEfDGCpmUvqKW6/vL7ZTL6+OiPk22NWbXGXW+4AesSuMPOLdaLtdQ0X3XYm60utyF7q+MXr
pfcuWQYomKcTYkttyD8vRvh5vbObia69W6Yn0KQb+VDRdXorBa+WsYoJRmfDB/rRSLY9TALugffR
bsDcPcm4iI2WI1OgVvh18UPZEPmCs+tvJvt5LKCFdbrjYc4/FEIxCEb6/dRz73Y9JGL3k8UyiErX
oPOkqJZWV0+0du/8ig6pISyNImVqVIAmo9sP1PXfHV2YZyJdWDzSuRhiHa6F6zdUBz6NHWbOdhkw
8vpypYrPBuYRtsEp/hmOZm2Xy03wsnM4+RGLXKNbGm1bAF7ixGEIIKX5cwrCUpsnNPMOWR6+zMr4
uJ4ez5sJ3nGvS7ctbbnJZJ4XTexmDoO9tOmnGrVeWkFHZowOYpklHaKUxuXTapsOt9AiPnMEMlxw
VG89JdzfC94JrUl2AWEqi0FiezNBABK4nTyJ1G//VKOlWGQdEvTnFJaGV9W5VtfrjquNWtuPIFof
cyCrjvgCS1mVNWm6pKKVcFjqTswczIhH7Z0x00vfLLMThVicof8Lw8mlg1JVqfJfJ19u1cnIy8mr
WOM6BEEInDCv6wuiQTjgFr9JDf/qJw7KtCBzbnDlpOSBh/SA/N0e3x8YA7cdvgyh3zJFyKSA70Uq
0fUnTU+iCi+xHSZYu88QgNgPOD+YyikHdx+ivhzWQeUdY2S1pIhpyq1351NFi2WfLCC94GlmbM8l
ZiIorB6lHG0xNAwMtUjF6Q9SoVDkqsV7FyktW4janL1stR/yqfNX8NpyvYNrltHcWOryqzBUYeWz
P/mhPec33idfhu6GZAmHJHJmpWbk8tCCUUeWXcafuFDw7x/SV/1tpEfXWbZIqyttTMCojJBVsM+d
NSBFdrbPuQQziIUuxk4faoyiS1V34sqjn3M9NWcRJvFC7RoywnrExwTjG5H5wno0UcZ7EhqKFnhg
VuWOEB5aMyEd/LEC19TjLBHL8g/tOx8YLoA4S5Dti53kc5MrsoEQGWkubhe1D0VQbUzb+zR6jHKh
HPZ78FM2x+1oRKp6swVlX6gREn2rj/bzriPAcACoiiWbmxkjR27CO6I2OwcQfYQWZDMfTu9/IWa4
gq2S1pLyj3oxExfJLQd5IEn+cxbNOZhqrtow8wdMCiNeNzeU75Pw86ZOVxD6PUqgPuMlABNnvKMY
ad6s/Zr5q4AznXx3bcypDou3LMkF6jvToyaSP96K9JTWXZx600+i1kNVtNeA+mDhef5GdIJmCllw
CactUiqDH7k4vdLiTmKArPhEOOYtwnfHhqF17LwUV0s4KjnHC9wslaGUxyWnn6TV1AaKVofZgUwX
jlEQCXUlo9QWGPMq8P7cSV3F792ShKgioAb36pYfHE0GRLkOZEhn2OL3ca/89RXOo/Hlc5jcru28
yr0xGBrCrtaZrIHgN1l4UDa947UferlPMElIQnY9e/V8Iwed2hIBtGBfIMjhadNWgv+xXjVHZKc4
Q9u5rQy72sHj5Ezhti2B4j6lZKs4obdCkOcgWrziy6XVipaAcSPVJYBIl9WZve9tVonN2446ED1v
Iqdss6em7cAq4PeKU5vWBB2C/I8PrBsD5U32EBehLaNrx8Qwp6ScOy/GC8N/XkkE+oRXl1Kj0PZh
CiXlE9SsktM3JkKoru7b9XZ/bRr2tzv+gwIJamcLDCDnJGggn46nNxJH2HUZDSzEa3LbbARZMfWn
j5s5s6WYY4xAL/h1BArR+6I/iz9OYaSNUrISUTfiCV6BuR0Pkcm7LReSgO6Zwfdl8lNRWbaha5mQ
/sevh7jx3YNNODunciJEJZNHzA4nHf+ZjAWzpCC8thcICakiP9b0XgtHlB2Rre5jsNJsKroMelfM
/041UkrmFr3MAZqXsaD92gJq7nu2EWRBSOEhd+ButwOBPz/S1vEJjnXQ0Y3YqoP6tmGjQ3TyMycY
35pLhJQlzpoNtpJ81ukJen1vPrquUV8U8yRHVMNroWccoqhTcye9lK1COEX2RapfyI5o7wSSNnTk
6teD8QyHX9GQOFJmDeGjblYwuxV1HYSttQUUebRltYVRTiiCTLhW7K033Jzcr873vbL+QDitj6RC
IWgDHKQyP0vam79QYBVAmGZs1cFwyYE0h68ltqwBtfWbB5t2QTZ2VGXe2sFRTy69642H3CDWfpOA
5heLoYuDH3xGW7yDf6XTvu3NeI/WRXgMB5CR/Lh/2wOe4L4rKH/mana9RAEeLS0XUv+4xu6p2gj4
FzbpWaGU9iOd8EmK80V/a7LUXaH4rPpyPYy9qAoIVstfrsJwNWcGzcLjPj8EYKNo+egKKnfPvAIn
JqlYt3MD3SqZUwi65Vk5Jo3pF6Uv0dkL8YF4mnmwR3VhxpO5BflKvHw0crQkIVAlEOinClbZojMv
RnzIGuhRcUxIJReyIwKXIL61DzQj1wyYj7jlt21O6791lzA2BifmpHfx5sNLu4SjA+vgsl6WjhaN
IUvS+NGBRky+tvqecy1K9j/sRN0gm7GpBhntoTmn36Ma6zPyWDuk3saw5prQcsRVlmwTNQFIojw+
CSbG3Wz9MQqItFLgDW0eWQdYHLCNeeAhEyYt2TYXmrnNf2pmdr9NqTvGVkazYu5+Q0ExKSeEVQxf
77Pw/73yPpVoUTC0mpku3i5zpii3Ba2yFzZ/1XU6Ql3Un6PdoUBxmgK8JAUIHTJ8aAghUAIlth9q
9d5iaBccL5gWmXvucAqmdiZfNXHvboiYZCTEsHUd4rd2dk3oprRaa+/oRMoD/FS6BJSMkcQ+fqTB
bku+DWyWtS0/+z7XRX2KmRCafVIuduO39aYgU/mzLkrLzYrlozUz2fA2FEhPDNPdLlE3tLL2zJs+
6QpNt+N63Rce1lLeYHOojNzMPSoOqaUjwOVFLn6RQCUmCGkzR9u84w57PQUZ/mqzUVXLIXGP8mGH
c5Zxuxsy+RWOEN5lKrzV8D+7v2y36b+yks/DYqcf3WAqMcLs2BncGJCv4lFxZRxrefWMuhzjDBAj
LNy2fRwYV2lZaAVujTgEfxGaF/gwhrF2+43IlA4IJGbw9TH+mc+htWxWab5TIWzPwz+zYi8L8Z2f
0Td3iNz3t6TuhW6WOGkZ6oEmrJuASjMyO0hOZ+9IQddrmCMo3dpT25VrUHBtyXB9aATMBIiHRDIn
FW/2Bk/R92S8DVrIzsqQR/OyKd0phRdgToxthhJTssALDpgRvzNC9xMjPiCKnR1/aoeV9jh3loEI
X7a706KuQ1tEo7jQRalCKG78x9WATrT7S+8G164D0LBLaM8t/u3rsThTDAD/w2ZOUt/6jcC5yrmk
kn+PRg4zOAquBscrILj2mt/y2WojH5AkMgAmMICdWItJzlCYR76LJTV6cayat3ea6njwGt9/MY6q
g7wZ20ThRQvZRIHwyb56vbDR1dkJ8WebBwpU2kGp0iV4CYPEQbbuJYCFpw5qZvlWTjPohPUY5n0i
hczfH1qCVyzGgatAqSsjOR/FfKjtGyiR0FYugU/9PNDBAPShJ4GqnFdh7bdMOPQaeOFCBuJIcQR4
XHEwuqT5+AvgBG8/Pm3ugFvBR/Ntyc1OpA1gKTJMlTe6I6OZoWxkOT8YIK3FNQaXdKX5ZarE1Cos
botnfeySlsmHHtEw9H3yCB0PV0pMvlkfzVtWtJ+o6A0J3Cx2bto5gzN0g25HhwxPnpj4YUS65o4o
N5Ru5nqJVt+P5/o1SenNwTToL9RphBHOiiBAu/NLpxwsH1bYGkAeRL3RaCg9LBtvETAaBO0oi0SX
5MVCnKAi6xn6P4tcWpaGa93VNnTfcekaTBBfc1rT8/nmK/QAsRG/Owed+r5GHaRiFU+05t8M95vO
6Ubs58nRF8nuvIJ2QemkgV809J1SoTadSGUyOwjd1Xi6GxwxxBXB6kQMZiQQOAuEGaDkVN4DPZ4J
rXzW8u/NQH5NLwJMGqbJ1eQ+fL/0uhcddxTbtl/NtxOy2yR7LSKHlHXIP/OXxLbxsvekBHNumTc0
ehEQi/XW9cRkhr6bS59s/jNbaF4ywFE+iY3PrOTJYw5u26PDOB+2zbY5v9eroSev7AlLr48D9V6m
6cPew/5IU3uJG1SrsgwsC9mOeMFie9k8/BNob7NSaPkN2g+Hp9J5FlLeg2RPDOtNgOFV8dpYO7UZ
qM/OW3MRJA6PCCmkQ5uM595jMFo0M5LBuC2uRh5wo72zmsJDxqidmDR0bFAi4Mhgiejcj0ovxSpc
ZKSbZCxUcxBOMqgKMvLdXXM7lVpeoT6OmQSDl7hxReHq8bBTFW9FxKqI8EchoCIz1esBHii1Ky3E
l4NEAl6A6RiRdEECVeBfE9I19hpKMMvftTy4PcwhzSkdG/8fLYq7AJZGnaa6CvHxgD4310O5zGq0
Q812nMJxXZ5tbjzg+HYaSza56UHBpXLLtTkYG3QupqzmEwhROrEBN1aaFgb1R45iS7MFF29B4NAz
3/mcWQxSWJQBU2Szn3gMhK62wRMx0fPYlL3kh4785dZqlZLU+WfUw1VDPfY1VJ7/yT3jK/OnGyxS
1l5ezwlO3/p2s21p8SyG29EfOmQCJQxl3E7P4K8bV5crWqu6rubeqiy/NFQTF6IfZSeLyG+RyqyZ
O39KE7OLqOzLGgSKq8oi3U++cIPnKBoCwE8oeeTmr8F5LtHRQTEQ2I2wyz3IBVQ9u2AxZ0MgAiqO
8HIEFlM6q7HbrVGwZqDHx4MEsbhRuLOH37at1z0EMEGRZd2ugBWF2k1QlY2bAkr7x6gTwZWQtFrR
15GaRBkd0hnpw3sstorBHwj28VmX0nuev9McPR1016YGLm0VjKv3IqGRC4C1sXDJGHG50GbA5SkJ
OECQmby2VAciEbGtnDw+GwgviGhf6/hrXrxpbf8xO5TMlfCVNHnzr/+ZtJEC9czsv3+j3sTqRLxi
/ns2/eJZqJWnmYYeglzwzZzG4AczrLFo/ABRR7BAbS0k8V/v3y1b+BgsWeEKVbfeF7PeOYiHxkLs
0XxnkPMnHuR16XnuTr75GpNbZzervloNHu7l3b0LETK09ZuN+ydLHoMIpx5+e8ZJ912xsAzjQ2d7
LC3LxzjoiWCcnZB467RFpnC87hcQGXbfue5gYxsn6m0RAujdG8uisyzUauhMjpTGja4jU5mCgwnz
Q0S7mq0+8XumFde5Yx5AYC06Ndfjdj83msQsr9eSRSvTtPvUtVXprY0MG/dfSZilxmrPNqOXXVE+
rvP7vfLtB7rw9gDP3+X2CkUI7m284WgJ6XvOvSoO0OiZ/uBRd82/LqTuJ5U4DKiGWq+buu5Xo+TS
idAeyzFh1rk/otE/lUOlDwpEE1LcSNi4SigliB4V54cNMkaRuzvZhENMVqGdJfqo9iO9kZ60pyI9
h0O6wAHvEYIo9CsKtJMMsihx8LXeGa6ExL+5mcPs6lJ+qKdZayFK35+QKB2igPZTVPdmHCsoTzvV
B667MGyS4wLv0xGSJVY4m7POuR7nAANhZM8/5vlGcOvUy3zqZwLPZA3EnbJS9voLKGryoOLY+HXZ
RHdcGmuGAPR78jp26NVDkI3eAe3JIgyqFpqVWY+OILWAu+xxEOGOAY6D3vd5naj/AkE64/VJmEDO
7NPh7KPMehFAlSaG1EAmN+PC57Q93pJ6J2V8mbylf9o0J4UAUTdPgXhtpVcQd5f3fsOT37IfXONV
NOEih+u7ndgKPhtmr4BVPdXLxQkkzdAxygOvPVGFnGw7ZzN4gvK7KACRwgSbBhon9Crjk9X+ocRe
cfWM/enHCwqg0ImDDObbn/bZ78O3pi/cdAV5i/fgnfsBZRVzAMPB+CsTEsK+s+962a/sNBV2i29g
UJzCTLw/pJTEwgJOrCEmUm1VftLDzUkWikwsvLohOzu3IfSGbP8Cz5+4UkJmVcN+HhFfXPlaeuVZ
SdPm7QYJ8AI1umOGlqDYzYexQoaGP0QW5/3WG71VxoldKh3RQA3wPVZ891H3feto83rWF5w2Nc9I
SFcvqubWm7LPggZdhHqg+H7NV0YOSouQLL8fck0GODYuTX4UHbNQrpYaTZ0eQJHb/XHSToB6YVCR
1hbMLRTUMKnA9vpTMKWhc5B3+8OpIztvnobasQ6rFJZaA36zYANoLb+OpaThFE4tCg3a6Z7B5Mmq
35imYJvK1dUw3rr5nYLEocnhyzwBzfJRkKM61DAcM5fBl2ogaGblwmWC0X+zQQxDYl/0ou015TLi
ewmWrLLh8kLVPoG3k6of2GSsFMAgZr3209kp0tFsgBLvStWhwmS5/7I+9M+7MIKHovA1OuSwlOZH
k6w+bf5mIX0PZEty4ZPcyOuP2AUt/lNqBgmQ0WF2obxhCsFzMkFof71+NRAzHYJjIdDbKlcfQG11
A5kXEmn6pV0ItmSvI4H1eP5sIV/3R+JJJ+xH+vq/rwpXV2Nj4KXleo6IYT/PkaiXfa6y3cxE43HD
HkKTtZy5CLBZbYs8rMHbgLbXHwAtVaiTAUUVKfR5yTTScmoWc4IshCrRe6qj4mQbNtxJr/jT9qak
yE46zRHBobRJD8VUkoQdvXll3fP9xCaEHCsbjVxCTKcUoSUcVWhycAPd+R+QZ6CS32DnnZwSC64p
tQNLypCZtxF6u1dkbohEQl31fx4MnJQ4z4nNaSVNGrNejal1JAwdddPvWm6frnIlf0cbaulFwmrM
tAqc1gUxEENMld9Ndn50ovrPFgO/THqKr3uQJHRlqTmPkySdXqU47iz1LefVixIUr47W4DyObEVN
UDbb3BAKQyzMwT4qTh5PpyBKgAORuv2MxfNgVnRnVf9fT41UMvEgg2DvxpnioXIxcQJ0eTkuc/5q
S/sFOiv8MTQ83FuQZP4mMfXiw40U/Bfn86i+4tPaYQyaiBc9OqPnSI7FHaBsydvwpBtc9XBwxEuX
hOb7UQrQRI1McBnLNS9poP+e+LQvVjKXHxmEz5yFeFEPch7bnISDldykFLI+rvaQsqk2BjtG9Ehi
XE4oVLLqGKef7dYyOaxa+QcuhfbKDfm1EXEHET5vfRP8l0+4kJkBEoc0ZfUUWt6IFKoFMWMEw0nT
tYQTMKcMW5kKiNbzLghn0CDXvycdg469JBRUHQCiwX0VsYSbDT0n9DjpuGvUVGvTxh7Zq5f/KlDd
Loh12J3DOb5cAthWO7axpwNUMOmISNl1u/CbhULi6rvPQRjZNMIcEl4KuPiQlbBG9wKr587wxSpA
g6FYjKwY3j7XfVZ41dyt1sH7Uncoj9ct7YoZS5UAUl8NqVLyRPgvVV2B4YBzXMebTxOfmXD0GJyZ
B2Y+w28gTVd5btbyeAivwn+77y1RjPvHrVZkEuSy2Xd/95wNwRVC/adicQE1lQ80JdYkgekkL1dr
631Qyu38JVvtPikUgBIaTzb7hKOpgQWPTQDngfQfIcLifUn3A6G8g0sscPjNT9fBqDmS+dbUSiEJ
4dxgDMS/c5u4GXQ05qsFpk0wdWw9+uIJmSdkvHXfb+bibRZ68sJHw6pr3BkFZHDE550xhVzwrchj
ByDcdBlEdzwfoBuWsBakgWFwkphalmvsBbs3naATZm4ckcEGXblmlk5KHu88oj9boF/wodixmlDJ
JfcpnOr4XgevCdCqyjworcUDO3HaDVib40teWhWCOx+sXDVyyz0blaI4R77uO5M15LRyNMITt2rM
Yw7xh/fh0w3lj4MAPcat6SrM+FU7GoFLfwa2HVZI/kgaFP11hwDj+BQUwPmCgw5Cvyj0sjQ2Iqvy
Kuw4aFpVotyElEGxeFj1m8ViAD7ycNdansX4kXQ0HDwCKwqZXteL+RW8YFWhTO2sCoal6uP3sPml
SuXOEGc/e7XdbiuGLJvQtCbwC5vX/OFTItqqlZewR0t3T+5zFswb02GShjcyfHpJHjlj9l4Tghb1
PMcllziskxXrAFUjvBYnHOsTEgGdr6rkwQkT4uHjuw/PpC45EghUsHf8Xa2Qu4nz18p5kLEdX1hl
UU4eEq/kXrkBC6V13bIboxS7pLtSXaen2sPHSNaLF+TMalcSsH4rLBVdBcG084PPxAGnTDnlLGEq
KjFY7r6+BFDFzH8mxN5029TeZJJfSv+ACcEm59jSFkJe83+vkX0djVT9xGyEJyaFekrS5Iq3lmgX
FqedtBAsN0UXPzw187hfmbHG9Fad1qzD6uYqlodocDcao4AorZSPG3bMloeRupdrXE6JPjQDK8W1
RNvagzBvE5mHuJwPdtBujODHh5RvnRflpmk0nkKenS41YAkZml7yhWfZH9kO+rDTtjwCRGpuRz5l
Qhtscb3BiQKqhN81JTetLX1jntfaFLCnUdJSO+Lzn/fINu5P4B1+x65Nkfa1eOavFacVC9ACffmC
1eYMsNyccYtDWKwJqsimU1aCv21SJCm2AsdUEdJv7WIJi+dJxPPt4CtMJMRZM8ZxLt7OuFOMN2oV
lRA1HnFEHDJ5Cris+dvbuKZGLxaKwN7d1OyKRXTIoFVfSfsUww0ypDmLm/HJMEIM7yfvo7OCHwql
ut3kblIW32EyVrOroPCczJ5uf/3wVcXeb3K6Q+mEzCJ80P+4x8my1WMgStjvNMyDSC12V/CX0h3I
GknQ06Fxjt1kEiPC5cST8hsjfLEPTeITZ6SVgXhDFwRooYowUgplA+8G58NsmpwHbvQFOKQRrUl6
2dWc7KwkvDRqfvl7MPb4yvWAFsvYJ2uzTznZekaWz8+5rEF699x/IODyFP6SJn7bA2GtQKETfX2c
I7ek4Bmtm13C8Xm8qO3iNW9pfndrJW6KseuMk8FvR4GOxFSMWu66uA3iuXhvsfSBKo8+CpT+TyRF
23+avC9Jy+YikBObXOjUmouRtAchSIVASXLTAno7gYqG/pk1mzX+fhmR56VFKMArMyZIGetc9qW/
Yn9d70E4L5wfa1tZxBWVmE1sHPdevbO6C+U2UkXewfRmrLEKfl7HTVdsZBy02njxFFBDL43SFAof
rXJxCfnxzXr3G/5xElqEra188hqGN4pse6ImEbFLjvLS/56rFyQk9Zz8EGsryT+DEp2J4Qi9lIPL
7FOD7pM9m0Cuk0OSG8O6z4EudbFWQnTMjkX7iHWBVpc5huY21mm7b8H3ceTMqaNgvcEoywG44X/d
PnEnw7NNIA+IH+vCBzDMBcEemqYtGBI/pJMEI2oC6LOt5tlc/Dm+oEZvGzHfzgy+pqkpfIPPefeg
tBdGJkcuSXhUuljHEYnjcvjH9A802RLTLarmCZMIaiXlLnFWOoYs5BNSQI36pGCLcxpx5lKfhCwn
2wnYp+rA82Gai0HZLZNn85qQqDevRErV5jswkbkL1qonL8TM+SdtiGsSmazspTjRg2z4whJRjh9j
ZllqGjqbfu3n89hO4pFBkXQWY213Qxs6nttHbITkgpcaZ0DN/rg4tRdB06lOPT2aakh57kftWM4B
vZvLwjC8UCduhD4d+FOqSm7qLrAP3LbSgRbeENjDBH7yn5uKN+TXSWbHGpcdV7pj82TTG5AdhMEA
yb1PlneEw7XeLzzE7paNYIp2f6mPdPhEb5JYqn05jChyjRCWrhZoFiAGOTgUANQJB4CcrpKCmYtq
oxtB2ghUixrXfBtZU0XWlgBneIJIZM3ZCQ6zUS6XFbkeU/DR4P/2L0NERBGFi5P69Dj5utdw+0Om
uVcXCnFx0fqmtH9Qg7m6m9KoNSSOznMGJKlTqLDdj+mKv2GHgYB8mjVcVCVylJ4fuzktTAILUwVx
T/Q9aNDigt1IOo8SYBJ2jpG5y0xkfitaeCBow19zSdO4YWyGz4bIYJQp7lGSlgzwcTJLaj30EXgy
hCZNC9Xfyyv2Szr6VN25t8zcvKR0WcToUVWIZsI9R8mFVjbpm5kFMHlkKGnBelWn0HQuCfs3wq9I
dxJsZl4mGwjU0V/KjcxCwEjwOaayT7QAALUJz6lJGm7l0TAWz/LpGeMO/QFbIOwS6959/qEnrsB/
Gx+1LdcV1iLQYBpnUX1Da1YIetemZqrit5RE4rP7zFw789Vj3mdZ+6QwVRLcx8hpE4eIkCJgQJ2W
uj6GnBoNnHl6o6MTZxTtPTYtllfwjGcKLNUu32/gtxVqGUWyS0kpYMc3RfN53QNHSqVPZqYehPfQ
aqUUZA+Wb+JElMgAnlgBTOxCIY5bbpS+A8cAI+e5TXne5KaBA8oRN6SrKTNaBDCLLhAMNZDUThn0
qpbDO+UimNETiJSlE8aZC3hx9o3zWJTGc+RO2cDPOEVwaPEEL3zo2HvzbL6PXZiKjdzsr71TFyb7
alFN3hHqTineeyKwgWMC32HXWZueVIibDSZllp1DeEEtSnamDL3o5q7ITB2izs6CJ/i2BavzlrM4
8hvyxYW5T6g7gdDMS7gewBt6PRKtQ6uDFaWLPk8KSqnGNsevbp2fC8LjgyzXsBUJeZoms3Va2zv/
8bGSFX7PgL0RLQMYELp0xoOwsX8yC6T7R7M9OI31gB8QPfN8TvZcZ5RBy2OieBgwxWIDl2RNc2Cg
uQn4CfFI5+doCAi2CwVVOIqD1B/7V67iakJ2yCVUxFF7FN616CwFaKO7sfB8Yp7RHFX9jdq9Ee6t
VuSe8rcEhJ1ScBaR92i2eu6xq/7TACRWUnkmGV2pF4Fb2KkUUom2niyuc9I6OHgQmowSRmDMJlSI
HztkziBT1gFKeJqNZT4A01H8zLyfVqmRz3QbSDnVJ+ByFK0golOp0H9f4Xmxu3FT13Twl1b1abEz
Yzbm8dmMJ94EaeqfF05n9kmfN01AtwxMql5aLs1OS9GQpe7LDjiGgpaBkAr8hhTtGbCY7zstwvs+
toRUjFOc29OQVmPJQpQxr0lyByalssfi5yCHEw2ng9OOyuiBHNC8O3gDEx8B0Ef2vQEUvYNDsbbJ
VNydNWJbHbi0qpQeeQ+lFwGBffMs2C0a67FiRvrzraTgiWN2wzvOdM+oo0SfhNq62mAKA7zOWB3U
TUZI+bdEc4vL190JZGvK+SkwaFVLNA7l3SkD8JycGi7LSa5x/fRY29r1/kRbHEVpbAfMHU+DunKB
lekLc5y0/3kc1wESi1x9HS5+6tpQDMDVWxZjZZs9sX3kodkgvNiipLpJ2KMc2lxTJMKZPQRlQu0C
76qOI4nlleWDByGMqfUIqULbYm0jM1xRTnxP5Nt/dFBCsvd+k86OLBlryN+1mhohRSRR6sQ9fGWf
eYN/hHF9hddGLO99P06tRh87pkgxmxp+U8WM/eltufPllFycI4ieGylZPjM5b86AqWcdjeCZJada
FNDKglQhNZY6y74NHj6AWsmHTH8sAy2kNZA/8F7+w0u8bUsxStMJX7oBLnvVQZX684RIBvKfYtcA
AESk0J5J7UeZMgYj4+9Vl2XKCG0c60QtMSVlNaLVlRkLgq2P5DDJJuGDASDRMrosBy0bm5YRpTxc
gNYzyDEaM+SRG1FY1p+OdT/AvNdNVJbEybpdYnR2/75cRQYsMPPTAOTSnn2YDjE8w1Lb4fTHendK
vLh7NgniyWVRR3ceryZ4CkCpymMIzsbxGmRqzLiz53QezUXkXU5nc13Dykb2V0G/D8VgjcUxlh28
pJxnWQdx7cK5m+BUXHKyVYATJtvFPAwUIVz83PquytvLiwgqFX66C5PHKfVev/p/UK+MtjXA3byy
WF9nQfmsWFmk3PMcYTiT2CBezyac3NSUVkp9tAArqM+ivVueHBjnjVuN84s7hsAGNsb7MvC+2SPm
jYd3e82klES0HWV4cTuEZFstrIbeKo/FjENOaLKF75t9Hwi+k/d77pM9t25OSQzVGd4GIO1kXtch
9Er/HhIeqfeJmvS2NGzgIxMd/PwARBeYlwCDZZ6Fz5I/5Kagma55Q0aU3PdELgHnzJ5DYALx/XWf
l2Xuz9Xm63MCTH5zY8owDYNBpELG1NCblY8LIcK7Ivs0K26296MDmJut4nm7IjyyMHuj+6/DbRp4
KVY8jf87uu4cNXkxlM6Gw23Z+ZbwG3S3P9tilyToJ8tsXshG705/JOj3Nu8dzRPDixuN9uskomo9
OPnYE480DBunXrRLR6YEh12z1+8FyATXmmyWtzd7K6vjh8AAhUagYdszVSsHXrpf4BMU+9p67wqg
iTodk3Pcrw9NLE0LloikDSR2lejmvk79qcz5Tx3jDjxeuy80xuzZAIKIlpVNSWt71D9gqd3Yu0A8
hL4eATNFUPpwuhiHIikFWhQpPVkYjzWuI85efGlcF0GtFKLD9Nvi+IX4cCL6hHaVaKLDuGjxXY/j
uYR8myNDUodh9blXu5Tbnnc/1NcOcUW5GtpYRGuuAARqdNB8CaZUk4KJOKXhsqZJMQw5Bm8uSKfy
NhZUHtEm3TKYVL95YPQ4TCK4d0gDok6FxM8qC6mz4NaUn+OtvbBjA3Zzyh/RLkuW7J0q+jcFMp1Y
Q66kmqI4h6PdLJPiinGEnAF1zaUrLypqxN1/AfthMZB4VsoXm8toODUKZYm8gBL4ogblZyU9QhxO
081hhVon8JlHlNzP3w/0XbyEoMp7vObCONeuH2Gej3pAiP9VRcYiNipWvuV1CLZEtOIU3Mr1qkQr
+XGRsNI5YJSxHFv25vF77wmkJuyJbEzV3tvvkfq+7r7aXNoJds7GjdZJstmflIk+rsiuge2D9X5d
eVRHLHAoKsxWMTYeqAEda5254FO9WCUrH3z4WxLBZ3IdhSqdSgEXBF1Ze3AGMzR4ae0dVZQwOULZ
TjlD7ZCKilufR2xZb9eUJXYX8RBAxHwXAd7MOUcdUkvQAazOnryBnkM23MeLzYlA4WlVk+e3AqrN
nd3cOU9XgBSeiQ5wU4CFXNtZ0eTZGC6qpBwI6QXr8/q4+SRDAnvXBLP0qnWJzoq6QrSQVmINsbLU
9s40ZxaWGfKYDByqUKGzoEARVAzVFbrNELXjO8LlpwoON9Z7WQzCqFyjXCs3GYxaMraSFxuXcnhd
qAJH9M0PheVXiHOHPEC+36siLPm6GRIZ2xLr9CA//dL14s4y/13id2Vc5ulPn/TPiwbEhiTeug4A
yPRNWLgeHDK1mBmILrh3hZbUvgw7VXvoVn8H1Xhrj5a6ATfnUx8zd586GllEj1YG6wNfaOjKYYS7
BZCvE9NG/o2WXCj9jgrHfmTN0GmmH9QSxDF6WfT3YzfmMhKBrhvgmK2BlmefSlyhNZfwvrY9JDoL
yC3brXkYYhSCr/aFt+5uQ2sNXfmwdtu/w5n1+ji2ZQgncnAHQl6dTl+v9WxSe/j/b1Ya7AO3YAoZ
ak+Pg3qNWrSId/uxdXS3qXCrjreSDhdKrxGYcBzZg6HU+qKIuKO9Y8vw1uGwS68jU1PXiV0dlKgQ
JEKByd8EfAM3bvFK6ZpknKaD1Uo8Z4MhTFSCLARj9TXyLv+O539WdwNfqw5S9ILrua9qTiLmGgDE
sb6VZs3OGjlGUAdMRZjNlnU3vXuBHuJLE9zivXDQ9nr0CHL1muv0YzsH26UWFDcQzgSwiJfLsdf3
hscy3dhlCufjt0aWyCUug+/W0XfVDNry+Xo4H6e47mI/lDYf6vwqLlUIUfPPJ2onP8UgVIZxbLJV
9L8rYkZNQRyZ1DE8Ed2rsT5Q0hIOvQ95U0aus5bbhywWtVZMp+wgPJcUv8fd2YRjW4z6QiqNqfPX
6JjylLv7QB7QfXVToGM7ryIVFZSLyWZKNKilUuzasF6lqK14tH5qJOekbzAkvJ3q81x77H3ryb2G
bDYK55X9fN/qADJlAA526WWb40Qw4+4yfipHorURlnfHWvtiuM7UYXn/ejVGNDjqW8TYldyYo9WR
VVpppBCxF33WDnq6ku6phxOQYpMuj45SupQBRciFQzHMXVhAfhQsKLtS8hA+QE6RZRMAMhSP9HSy
uiERoWFKtGz2krZt2MOZuz57P1LYwEzhIHEqZ1x6jGKB3IMYrPqWZgnxCeNItcnb/9oIgMTQ+7YE
9/ZBLiYnyAE3jwx5ND2F0oN9bHI3PpDtcW0UZUdNUk75F7mO5xtL8BdMrUDnKKvOyPde1lTMp5Io
4SPf4MxK/WtiTiEXm4HwCoxr3hchMH2jy8RyRQ8fF+YFVSgJ6P6WEAByCoz6fCYPcQCv4g/AtKLH
R/9PII6cnCvpgGcGK+agOhiZW9Rd7yq3cBqGa1EGUb2hZNiaZQqbRaobLsoklFW01X5B40r4/50Y
iDjsZfZMvb1FB4I1xxSTZA7Fg+Zby0s+5aTaxC/gHBuyQMZak1r3ch60ADROnpTgWR0YhU9rnt0z
tPfjtcn16e/TRCZwfaOsgGV5TfDxg/qcG9YEKI0wgntSe27M0P7u6Q7bVyiqgBGMm9wzIHSgj1D3
BeE9QhPD/cCvoR4NUheotg4sDW8XutdWv6L5y9ho92Opewk3roT560W7pqwfanNTbPRjaOkxMiVQ
liuYCbLdkIfzbmWALbAHr07Nltqp8H9X4a7AowwEyuaPWNAt5JukwH5Qw75jjrE2D09BnlrFfWrG
Eu7HO3C/ckZ9fkT711SQssL/Xj8hlrM8fTs7NC/xQ0EfFuVS68kNrZBiiqgWCSYYYmrfePvqpYls
N7ujGKyySrnO9kTyJeYYcdHFum1bet5vJVqnD0/0XTz2+i9T+p5cAIaKG/wLjxUYrfxFchyzPkoq
ydECB72hcpAjBIQ5+9+T87Urug8rTYaTfT9a96q0k69u+lnhwB6xBlehwiBNekzvLkZs+lOKsKen
06dcJq6yxFL2LDtZosF10bJ4Od3Tjd0YXlOVuTd9sBoW20vaARRgjqKabje50KVdPWT1h14ALvCn
BBLWSbK98sy5boAssHZhZWFTPgPztSMxC1NnQAydX1YEz4MdWmKNEgLxfAD/DxdbZFc+lTMORB6L
VC9PL3ElK17Uxx1fNRHgj6BgEGtHZ4AxM80Aipy0adyAjIaDZHrk9mOS9t5n2SwbNDhBKd/zFTIu
gRj1ieES0LBS6IzM9GzyqbQ0DJEzmqL83cCEdV3bpwflK8arG8G9qQ3wV5tqgERy6EmedBQaT6wZ
kBFs/ANIUK8bAoCs5pJhYeWn8owZt1PRZbFOQMR3L8pG995S+CvyzsuY+ecpX+pO8dMK0XKE6NJx
bvWMpkblsNqnEzAfrm6yBjVoSIXP0BAhHFmrWGQ0tZ93sFIATmIlUq1hTATCGqE3jTWc/cHD8VeT
7HZrajzTofcPLDq7t9zJLhPgBGF1HotZaANRU0kZvB69X2gaQOhSzcW7ubofdOYEAVRXyCTG0mSL
blf2GLByVNbK3o5gjaP2oAqJSfQc7nGSPVL9kWhB/0SaX116HVsnkvcuH3Jd1pm/1rYqqb9KytGQ
0nbigI+u1gz6FtuHwSC5dL08uTMXMn2PtBDcs7dWQIHL/Wa9NtN7QcLNI35HqCyhZalyb/tFbKA6
QnwuPE8yJX2FY1jmWwK60r/vEaIitPNociFimRxJQ86cDw6cbsRwP/gHWWg+tJYU7592gQwOi1mR
VUaaxk7ssdpfG8XQeSwiDe1rFqva93bsuzppXyx2KSaxREY0dJXCdwif/IsJJmOtD7WPhCRKplz/
aYQNmNkZ62JBSu83wdMTW1/4cN9A42HIDNuH9EmaqRVUGrThw9f+psX16mckYYIeN1Uzllvgqbnn
zHWt4fPB3ekIQuof2xFF+Jo5cUsxMJTiPdRux9+20arjsMdjMfzjA6SjuqiXKXk9/LEPTPfJuCVb
KKBBQdVv7g0qYKe8HRd/J0yL9T2HN7XF7hn3YMKRA6ud7UqCJF0QqvyZgGJDgBlOwex9mgaA/8Q2
KEkhVG/nVSwfb1KuVeB4Cl1v/09KFe3OEKFFXytTyXfV2YcCYhcJ5ieUDBWQpQQXYo389J+wdEhr
RiNV7Z4sTZYSMowNm2az54ccQw3ZXAqjCfEr9FolSEqW5tkih42B6UMVOfBV+2KqHeNo90QlNUIh
dMeeqqoB5eFr2z8skGaWOP7vIvCbf4VrtaJPZjhBZDTPtCHMyfctmVavqOH1uZr5APpMvP+IwnJ7
V/h2LLlMZH7dZ6BKBmAkRulweE4/wRbLVLmeviLf5cuNPd0r/kF4VPJE0HFTCYzFmPdZWNbNpMd0
0Y6nLGByJ93TtDwT6ctHbIqjjGfjBN8RBOld3fGrhfsC/YAOnl8MNVYKwxq4cCLx30lPkMEhNe4T
Y0xfbWkZ/dN00L57+kYEBSGuHPOLr5I3KWTadTqKjOdPbuPNcjKydxuzHY9PCO1XjXv+3sB364lK
g3FjSujSzV9EEBeeLriP67AiwGq8RwvT88P/vykAdFgdVIeahRR/0erCdSwJlyWeX4BCZniZvjLK
arGWQTR0UfUPAYVBdkgFJzekh08uQsPNwkyZ1NiRwoZzcoKlaWO2TH/r7v8Abkgeb2FWKO1TqvHs
0l/6N/3o0RYz8zM1QLG+34uqxJAuKZMNqfDnDdLQ6NHFfVGnXO+mk4zJf1YvQLtShVF7RkH8fH3r
BMbG2GKf9Xi7ZIO1WLD0Sw4GQijDS4BYsux8oHRWLCnq1k9BC8cMAa6qrTziJa1wHMrxUBy9Us38
rxcdSxIyz/KtXwzV8d0GV3ysBlxKAwyyaPFPvNMXWDasEBJcEp0pzA3wCbFangC49ZNpeifNVwsN
oY8I7FzPdT8mLaxFBxAMONBiuo9TVjYAdWmYAgzoEqxaOIsuqtl+B5ppjwoY+fY06Uk/cLGOLjPa
JZEkkgEGH2dIk6IkazkBoBL2GTbo7/6QM/3bw9fjihh98gC9PofasuQLlpK+k6GOi05oF2aWIgfE
ZpZim/YkqkSkHQATrI6oj8yhMOy8HgYpxvLlnYjlr8bAjnT1i6bmDrBOGehC+UXNHtA1T3i4kut2
QveZhw9/qcVjepdVjAm6Wgqt6A42ifKyovCng3VTCTaV0x/ZhX5irlbhfXwDkdK4jHQFgYMmUCWV
e2WpFlHUopNrvAuo9EupZxIv+CxRyl1WwXHY7YkLvV4J9St/3VCHTDCu+j+a87rQvJ9ismV/g1gM
n4Z0B2zScAzM5XB0lLXLcvHXHxJqVZDXY8A+87RQmysooasyRJd1iDi85MuR6v3GESRntXyKV753
w0GB6+Hf7wlO89FWZ4wNzEsr/OdX7h49V2E6hhd/Mcm+fX43+Sr4A3jRl1pguiJZUSbivdg5OREW
i+xWWi7swwTH2ekC8886BEnhLibhjAtc9w6OrP8npkKsaOHFdZ6REdlwsnxNkGTjqYnzBT382xPV
a0kn0lAIBfyedPj4Z0TgaxPvGfyQQng6xQC2EldFk5okoPz5xq/Lmd7Kpudp7uW8TKZKAcSlvfiC
tZ+0RR8exl/uc/XAFkdkk5nGFFpssUuslwxEIFmfmkburkzP/0H9guttAias3V+v/Gy3qnycS9hM
1FH9i0t1eMbxvs2L12P0raJA1P7mgcwUuqZ3eQ9dsat3D1idUKWB3xMjsMFad9qybsFEql4MdKF7
j9Gz5EOQRvHN/Zvdzv6od3vgtRKVysfghvpjTNEJS3PnZLudLsvfA1Qc1bPWG81Dj57TcVq10cxY
HTmx7JkR/ssW3FyQzMHHcrjU/X1+MmWqmGlUdFgz/mbMe+jScCTgJzblCiCEOi7XpOCaztsb1U9v
aA1Ziv2/sH3esRTIipx4+cG2uJM1TwTfO9YwvzZsJAZbRVTVhRVYfNs2kAtvS8ZRqr5qPkcLjh+u
UHoe3EGnwbYwIIjcgbo28eruUnYvSW73vG/UdOdvWUu/xFVBfkGCBu0xaeSs+hySTvXWIUaCJ6kn
SDLzH9+7PWQ4fxVwMj4sCrxtGh9QpEceXddpMCg1loun1nkdg8JNzGwtI1QvynHtRU6kXBHVdZSR
fr22lTRhI4v7czcSrxP8S0CvR8ThnJko47CfSSK5TQemtB1ekyOdySD4HVwCvEDsyH88BW+A7G0t
JomRUwtqq1757EoZTGeVSw4pLwYT1q9t2cHkKz7QDDXIur0ubUZMRcPJJsHTbhA4yjUlkdt0P5sM
2ghVjwJ5QUZ7ywxoQki+Isd53dctetqjrTY6iheckSLZSoAIQIq+j0Mi8V3ZsaBwMjErNKK6qgLC
SeqlxaMmwgNFnmMCGfu53hK4w3RyVn5DoQ5TROlsNPtvk9Risw+WK1VmJgMdJCvmW72oT2ODHPX8
C/tA5T8eY95nwl4OlEHGx29Alx1qiMSRmxnmxLZvxoZj9b84KrqeUcQTU3aCWU2cc0Ah+XZO4kpK
AK1UV8tArA7/JSReQz5EESJf3N3ct1Kigm6GuEtdwSieiZTW0KSSQrxEAdGl5u49LQWSZpE5ynPw
ui5joYkWqzEl9frKtV11OJKrxc6M/KoJi1caS4bfCOtnU63iyHUlTCjy/s7+7IvK/BsemD4Fo6em
EiXWk1xMLK1hvpKHD/lCHJsMJDew6yPMXpiOyhTQjtiSpLTEy8sYK/n187yOBwAOxDfM2vnaJgaj
peJWpMES/B36XmEnV4jcHZ/fjD57d6684R7Sk+ybActYaxeVTADjtC0290X36nwn4Bmn0J+h84ub
7ikebe22w7xdZLeR+rheZzh6Toqz5oPNiYXZI37wi3k1V9hKzNEg84QwJnIzQL3X18LoY0TRaYNe
EyuYRsKMNr5xq9pc3XFFfSGCmx/H53+5SyGCAtL89bLyjdueCZdfu9sb6rD52sCb6Nndq6lMSOoD
7BdZKnFQj/KbZoDrMvASAeVUOlLXpPMrHg3bveN/DMF4lt8jMuh7LVkDBBC3Qs9GOUABJ8ClYDeQ
Gtg3ltW48/RYyP/hJbK+b14j8cLtddHTg+ov1VoICm3ka6O3pU3eWOKGnwKpJLsAxmvWB4GL59QS
xtRGg7UfwqhjPncR5WHbZPthjN1HRBJAGt4TKNfHMusFa95abjLZYnBh/rUKJsqyhX7F/bKgOv99
RlhDzGpXjTv26wpW5B2CiaxcKxoiURLm5djY+9QsxMx835OFv4QuvaHozAyTxrg82O45CJIxDTEj
itDYfn/HTAN59C/SQMmsUdGe9TmoVGIkHfTPvfj5q1ea7bV5tWIzpNtdbB5iejSEE9z+LMw6+wzv
z3h5/XVJ/oLeyzHXYWQOeZpFDfAkTogLvQIYKRfTU6IXIfmUn1nu9dsJsWnikLJjXhWC+H0pDUsB
chwvGkIsc26rneMAA52q7IBSOiNK9gSHDAwRUjeQtXzqK5Ev9N8ZBJlhcB3uciiXCle9MP5tIupj
HsTy40tUrS8wm6GhifEDcVdORoXyRYAKr2wjNC1Sgi4avwXOsfjD5HKbsUYOIHp454BA5ehoSkhY
6NYygsJQGD4titSb18FJ0ZNgPR4OfGk+4N59e6kBAsi50qY0y6bQoKXVqbv7ifz8uHOcYKWy4Ssx
8qaxkDKn6CC9EkYHbvvmU7/WtR7WNMTgv0CgkHS2NaNVeOyQ5vL1n5bGPFWFbIzKYvVpXiKsMctu
Hl3hUiNZtp3MomugkCtXMudm3zaW6blBpqjAqULwLu7ixlblgZ3x34of7R8WzX4hPmYKpUBWL6+O
6snnUeotcBBy4xy37OLPBkgDyWVPE97vVZI9nZB0UAzeP9z+zVxSUfA4K3Leia+xOKDx+nPM9OGP
qk4URpzs11ECXibpz0r50+I9HQopzTHMGJYqipvTVe1toPww6MgBJ0zgk/U9QqrEo/DyoNcPvlkt
x5zpTtTGdThiMeYhG2l/QrcOaXGLbHWZhTEQyjMeQm3tliuqxAeHgALHDI6q8J4lBwU1ga13Xfrg
3GIK+22BCCz77YLvZv698ZC0Pdfug9hbKRKA8x3QlNS+XfrTbrS3Yye5jWViiKoO1WF7g327r8cS
6pknyNRd4DZWyKc1KHsr/e8p+oWj/efA7WGmShpGaT/UabN9AlcmGDhDfUHM+/emYForjtKTBQwR
SFS/INsDt8EYPwSRg36I15fsT2rSohLM6S10dqIuJQYFhKHfQUt7auFUZP7lJnm87NXKotpuBwKf
/F56bu2YRpaDvMQRJ/QUR05U1dbTj/MrRjz6QKuG4UjE9FjMCLyVnuDoEtbcekSR/2g9KnY6+6Ap
b6+FrGgL1Kz5vFF9Q8CdemBy8NNmjXemztaF0D2deFK6ttzXnCrNtrYopULrawptqRPxcM7vyvav
UF262CSDNn9WwGD9eAlegPvhepjgqkWnsEGJLhJjtA2o55dbkcWTADg5TGWdUd3tStwWrU28Pg7X
SEynvfHOhsfCjSMH3KeXAfliF83UJQmkwZTtwds5ZKd+2QeclW/OjA4xznbqxhvIoC5yhvIqFOTw
92sDEMPLZB7vSe8iNcPyqPDUIBLuE/kXa7HlzoNyekBXLU6MVuCVNirZya9F+pMvwC0SCrZLGLF8
SkoofwEapw/X51o56hk0BUxOcF4ZEuzML9dx2cK4Ypj4jWLf/teAZJ8hpU+7rbg6MYgfRqtXJyrf
sPvfARkHgjS7sr/6yEtq60UPqzhIxfbAKj/L9eRg2TkMoJUViycvA0W92/oP22nQ8KNAMgIxTl2c
OIJFhs8BbrTtk3++2tPEMCumT1hsjvf27zNrqqLcfg3VJTKp9iGO+gYaDkJ7lniaLrglFaXHKo6x
2cbv3ETD+LqtTLOegmuRUmiDOdsTRhg0J0VXE07NDsOk/BtMYqWET8Md1NO+yiwg94u4Y/9xBg+5
5sf5wikrZRujTCH6SX/syY2kcLjrK8EU1NDkWd04ou0dqXviNIVAcjB06tzCUhm7k3Tgb1MqTbUd
xfByxXhkwYJbf5Wa+Je73FOosp+A5bastxUCpBCkUmPepZsFFPGzVCkBQeNotrp1+HEHwBo3b7ua
omSHeQWqVGq+8msRZG5BZI6DEq4qK3po9XMIYbbn8SqhXVjV/iRIS2UTPmXGDEOXI9NARc1ZaNaZ
LG7sOUqmO9woLlyzy4yHmh0Rcw6YjhFamwx64NqBKMLyTnPUugGwpoFmq4fIlfGHtytpP5MbQGNf
vU64CkpmY7a3xbzEcJ24MxkLkIziDf6PM1TzOgcOPW1YhCb80LqCnZdqPstGv+JzAYdiWaIvXmzf
yZlJZlIaPNv6XnJKehcWAZFxcLpV20rl9jotMEP8HnR0xngKkyqpdvYnZvixiA6WZ4FALE56UO/3
h3CRYT9RKh5VMzZOVDrROebWFuKwiZE1DXQvS8tCSWBI9mrPIz7AiRIrj3N9zKaTOsGlulKS+bXj
waMt72BQX5Q2D53phiPitQRIui+IlFtCcf/HX4jYVPMUZWw8sYFGmQTvzLkmF26O54CPxvR+pKZF
YqUPsJBOub8QgHA7woIk+y12xjkjqiqwYK71fybkN4t5f7S8JMnjhsl8jesv5PVKp3XeYjY+w6pp
mSoXYoxtPtxpI0nnWtM70nBHc7wzKjXgYiQh3JdEkxb3ROir1Mwicf8wFT660Kyx9lQPVqFEhLfV
mlm2hvYTcbjADgnF3UiIoSJsoY1hYz5Hmc5lf8PvggMkYg3XpEiFQ3VGozE86z/95nVv2XeaI3ax
GcQbtelol+RZY8pEhJiwZYiITO4lhxdWG6OsjivA4b75l0Rw0oATjLX81pC/S+HrVPlQWTUMyjgB
ylPcgQ4elmU66ndpzmVhNZNntgOrf3GRCnEzgPbZjn7nc7qcniPt94Fngm9hGGgtZHu1j/If9HIo
bCxEurUr1ojYkbvVfNGjIb/TOmHTNp7hKOOyMJhYxU0OJTU1a89offt/jptAz9TU8KEhpWdCF5Oo
BV4Gg/5cwtKhNEKU04+JtkgBLIXJLFiQzajZir/uRUpsFsEFEVdZOTanlYTXZGTOgJshNxsBCtk+
xyhsRYM9ZqcFPDjtmobN1v/OnhaSO6PuHU0WN51XP2MyyMP6fuIieQCpdGuR8SG5mhF8TD5sAPNp
uij46FwW56tOVD8FfOL7qq0pwLnbDORbMgADeSf/sALZjsGAY2GpFRYylmo7BeeUzpS/yV1W5U1D
gRgsItb9QASCp/6wzL5cmOSQUFoK0nc3wkP0oAelio/chAqjEeaejGabcotrno51Ld0fx0ooh0Ht
t1mNUF5/d3r0uIBCtRMoOf2/4+CljdeSkhbmLG3E5SYY5cEe4K2x1r8KNZvGMiKR5JvuwHgmb7er
Po3orD1qeGqzPvGug4cY8oqoFBy38hg3GRQgsAas0kT5Ab5TuG81KHeDWwdPGeC+hpis+TKI63Nd
oiVXQYelcv16b5dXVF9A8bS/5LWVxafmJy+1eZbjQIFxYK3SbQsz/3Mp/2robCTg1E5iHPWWCmP2
FyITw8GxFPK7OPnFEoQXYqcFLGKaiapZcn2fiC4rVxzWU4Gua09ZHi8R65PZMsSg00MDltdYnaMB
XVe5sps2LmuiefQ6iS9kUjomJc6j9j6lBFSP2BVRLJn58kJkaeFzgFUYDZHos8zyw1TYcxu1xvRQ
h7fwKRWuqzJwJo07rUtZLrgepfwBOdKzgQVMg4DKkaWRizpTdOiHEk3K6rGVFNWh8iqQX5RmpKHL
wtbnKXeMF/eEFZMJYEx5a/3VP7u9SaEId7ZM4d4LOqzYzn2K3IR0U+m7kC63yUWcX32yIdBj2t8X
Cbqw5GcWNe/jT4WEQW114u71Du8BL/V/Ee8NJZxpO3g9flkktEYqvfVvpxJ/PphFgqI3ZRI9u2CP
i9m1FcD6qSWk6oERmpqrjkOkryJ2BniSr6bGtyQ2uAlu+/G7k8Scmp0Q3UZ6WI+CbnaGSEyIHa7S
udabe0TDF5M1bo85aCFi64QG7SwB46Y2eBixVKMQhIC9OTeLtfTVaOSOhk90GHjufvi5GqUjY47G
QInR81HMwhj4jW3mzgr3M8PA0yhoPhkLGuZFSNlNGBbO33IfCcnO1Jszc1Vfgpyuojxe5qf/Tyly
pQpgz1M0dYgDMxgIAaMBloV9VElzRIYO2a/UpfpIIw0si5wdGucQQW0py5NJ3Uj7uEJBPwBdqDW/
IswH5ZeZNJjPcUdwF63aYdOTI1TapAaLnEkLguwX16dbrTMkP0bwySLtE9z3+5uFkUFWMKKqhJuF
i2m3kIqrShJM39fqtdpl03S9I6VAlmohMghe84swh+vwTIzAmpHbHt0/mHzG/nipBZyasSqE01Mj
ybKhybEI90cTicAL4yxOctEv48VfUdHJ1ioONb8Ho/hwqA0sji2gIz6RGubBDbeSvG8jOKcyqICl
owG53wlhuWaHmwDU25Y/ft2qomK/XrI+m+7Lcowiuh7Nh0y3DRliqoqKZF20vMTIWvG1p8ZgcIBp
Pj1AgxDuX2LnP5MQX37m2RtAqquoAjuBYqDTL1vWR8OXUOU+0MvqVPTVx1nx1X++cpcUrjKFRBEC
D7/u7o7J0cEfuG441Ws53GwyCzWeaCnMDXeXc3TpewUm69+palI58xFjUr2ebOq8rQnPQTrBMUAl
OZB3naa0OtInPymRXjLdLpCdeUiSmiI/kF7Mq+BlttqkWzpinrcZoe/DTSqFKy4ykSrGEjd1P7Yu
eDwwh+kKqIj0Buk8DXidtH3WDv04hZK35T4v5l/5kxnpdqjlulZmqJirVkZzNoQHAuIrdEwanWA4
gsQzh608gTSrI8y56X2n3fYrCNn5eCPQnFjILYuNHVxP30VrZhI+fIUFPwSnRCIVCRfWFYBsv4E7
DH52ei8sQBPz4jcQGHGhsEVxQMO0Kf9KjKw9hJR+PSTS1DninfrotbDOYKqRB4NN4MPwQgHLCNiC
ytFr8jmKiPdSRC6CINsaUqLvEodga3iAJByHuQ40X5FiJRKb2bXoK00bwxg5B+EuUJIe1MsoIsyo
Jr6aNqVZt/JjIDjb6DWfRkAcA+YL+VSD4UG20GhwWyRzk1+vkSVAoNE32THCwvLZqTwyCtNeRM/J
/V6AKALxH7z6JspGbZW+fbbnnbrBwqeTFa1zbLG1w4ElZc6TySawlW77m3MD3atLN34KODzZlGDC
qjRsmV0KWmVF9zET6LA9ZDqUlJ4XL9QysckTSHWHDOUc9Ug4GPmVRmVYwlmT7EA6xBFl0AEQf3Ci
NG/yNCNfu3/zLAbxjiQ2jGClKYolgCGzZ3UTNdnU+6VWl+raMDQ2O4f+U1q3Gu/jVy3KCI/W36uJ
nXQKSCzix4liJLQEOGNmx2dI/M1VfSdB+PTF9kb0zFzJFSep9pc02IqSVD887gAmh/WROIPpdDBp
/DHc/MeArEVliVVaE4ozllVAtKzgc/L31wmstj75OEaMWtd0yj6mYlmu78zjjymSMRwlhTFUbyhJ
IDTYJXeJzq40Ts4CDe/aG0aFjfXQsyPD7qp5EwSG3Klezw+oyNb7+zxLiDOuCTh3EKwcMi7XsxBw
14f3+J6q12TchTz0yYRDDZ2vcZOtuek7PTX55uGnFRf8AesHLga+CkZ1nfgsqnTxykqKrFzUXkv0
jY+4eQriyCiIA+u1cExIK2IRyfD/5rPZ1r7sEbWmSn+oAcN9GY5wUVTOtUHwgjfxjnjdqfXE3ZEK
CNC0+CjjqoOGVuUb19Bs+KrTCuAgcXo1lT2HeOx+QXTwgfTeylGDkv7wJyI/coxwieprCVt2y33O
SU1+xZzWXTgfpW3su+2ph6Ke2edhDlWhmvl953U3AX/F5ExXT7litGWpSBeKqbQOWbCOZfx6T3h8
FeVkprcslrZDSn+o+RIcfUDxhZUy54dFJe+p6CEc258gLhHdQz4QDfmUF0Wclg+poYuVySDdLNm3
ukeEi31M7VkpXZyRfcWqrvJVRKNg8w81JRTSII4ZAJTnvPDB0rNuYih9oaORCc78IxkfWl5N7Aqn
ol72XAJGSLMoFjZuzlWQZ5yEE13KXqBx/BfpvJQnJCBpH59pi4G95FWzS+cqIvBhDan+48QkJFMn
j5lVIFQY9B6tgejQgrN/dy/uP4+aWQD8IfopEwAt8ugJgKViRv/NN5qaGdguyXVojGrYU0VTXACH
qcSXUwJIGW/cLfrQUd1aTnXqr/rWVJOeLT2c8+aLZrhk+Cn3WwUFfNrNxUIkXjBGrYwOCiJkFJdX
wP43cV2gbsnmGQNjznq/BDhcmS/TpeQ9MfPjgFXuaYr52OLs+vArPhacZwvaXq8KsSUlYplLEdNx
4iW7raYBxie4PkM4GK6LwqbpPXN7uHo4kxdJW5WC9hh5BfTwDrcQC8TseJENTPh/aoBDTcNDBLOC
wWshf/V2ZBJGxrcdtQBvSRyAWLwkbEyncm46d4TgG34RXzIHT1j8XyFxvNv4MLGoMqB9hi2CjNGK
gbWhzjh8HaWPALoADaCYX1jqoJKYXsghjotvfsch/mrofwOz26+EuiMmN7kuVpZH2Uc8WRP0iW13
Pj763cndvx6Ag9HKgWfv4icT57vDvGUMEcuOcj6SVpmaqoQQ33VCUC70nk2XmEOc0o5UE8g+O33Z
1Zo42bN1e1c1Yuz4YgKg8c3zXOTgAMipatMfVEzj/kNy2nX2fijOc4nNLvubBUcar4tUaQ9oDKro
OdQ9zwBv/Vh7suFuE9Wm/1+WvvXE4nwBO8e0u/xV+TnS1NR1pufHy9uaOg0ysuuN06EFds5P9RQz
++FAaXsS6tANEnHVWqDL1k4QI0V2AzyVQqi27CU05gsmXbcKvHwwZK00IYzyy+m1Zt/1sM0awVzy
5QFnj8pLpyMCXspuN/AG/Uzu0BM38zFjcctBZFC6l4ib/+EN2r6/v80ujYpkS8pUF1KB+9KQxdzw
BWnmJ/646HHdJaOYJgPdRcZPRfNksoWv1iZzIzpSDL2IQS/gfmVQAzgyEmDb+pmnKWRv6U0Vp6BY
ZGSgxm1E8ZXvtdp1m1ZAKKEDTT+EkAPfDoBOBB6V1I41nule1Vwdulphm5eCx36I56A00skjM4/o
cmm1pqcqpQFRzsL3z6C6SWTfXaB9ADPDPvKU4J2b0eU0z5fXHr4aV75YENiGo1TO52evvVZI+SJ7
xY1UAteATU5GRRDup6PMGhf8mFn/PsfblhfFAURIDmyrB7VCrDVj6TlD5w8cJDYz75HaqqSvyZLW
Krks19QfIdEtmCzcRdVjqPvVIbMSwF/nYamDbyJlV4gFMgQgd2msqdQCyMujtrnxtajF8UyU2awT
/FhfA8uWiOnkqKiJmg2QaRq+5lChsUBUAUaV3cDEhEsfvjxMf3s+fWOHcpZZKTlbqoW/9+8f2nl7
IKhN9r/XLA6l5gQheb9loNuTQ/U7fkN6v5qNCvUPDhNd434aF9cUGPm2vjUUtuZnB2Wpt7xUgtrx
v8sTNIZLEI/sPKEJs7rDbwSXpqq0/ouTaAHbpMFJvERkx1WtWhRPU6bNFwpD7XlT1e//jjpzc1qR
BWFqMJi7nf+cyHr6+egkDoEPYKz3WIObyXyocAfJCHjr4aKxw2ZNETvzVejnHQr+OUFC9BXyMybW
EORMggG7QPtVWp4XYP125wktcFtewHrzfTeujJ2Gd2ZviEslWQwWJT4U3SxQF00gicKEg9IRIrfC
uNpahxmcoakXShMp2HXwr9VuCEsJSmYsm8LvzmJ0aZ7V2IdTwC8Go+Eu8XvpYxCSELcr0zFhM2wl
G3w0PUJWIthUPLtucs8JR5qx7Q9F6BFdj1idyx/sw2FR5Z0CluLnUMOHMYpX4o+nk6aNf1SSt4pp
4brLXd0kF0tXF2wJWo31vpVRtOwYxkEWJhSj9jTbjKV+vHGWyx5rRA5+F1kGMWmkqnwmJlydizLP
I8/pXSkiyXxw/NXnlZCrsF53Fa4+8k9/Sg+8b5+OqHTB/SLxGf5GJMSDGL+ScuKdY5ZvMgU67EEO
pk03O0/NrPYy0Z8x8MjYFNjI5PPLylPCPVzkaW4+MyWZ3EA3ZPysaGdCkHdV7VIBcUXMB/VIUKrm
4rXZFZZP0rFaOAzGWJ1qrOopiLFN9cPT5qqYCN20RzHnRzK/KfpEjeIZdh4YUN16gAdE5VZPr6MT
tYejHe0Yid69+j3vUrL9o4EeyqjJQ48ZODN9Wxyu9FE74ceRR2qNF7gGFFMn4vvTZt9kphzsEhvU
SkimHxucTyXqqTfZEsfep3r0IAwwBWfVbVy6jwryv8nhs3On/2HYmjKQ1dqnMnrBMXFjmQL5WNNK
7xTEXdzTilBmcU6WGQLT4hczmtHX1zzQ7f1Q9K+KMRM8G4HWkrFcSpNbVliakhKxobIiG0mvur5H
N9ahTDNPdNExtsd//NayaQQ5hi37AZfUQ9hEVUuAAVzH2aDN11zrY82Sc8NQQPkXBBcrWSKZXnTS
PHS/6+HFoJuYdQBjTFilrU1zxGO2vDuRknfGpXQ3daf13cRGBD+1IyF5oSoCX6TjS6LADy/psjP0
pPi7HyEAAzSUR7O5YJMXoCxkHkbqevG/tANGSzoQhoYffzrgE9LgYu0zT0h7YNenCtP2JsEu5ANe
oI4VU3OD2V7AZd7VMUmHb6wPgUVjen0YD8ztlPKVz2JeNOxU1jK79bewL4a41AcZkMVwUbM+mRM7
H/kac0kjRvRY2KJa24XdI1ga7QSbfs9yIIXxWSTrSzZRAnnkiTHuyHtkv1hbzkF0YlHeXbd+hnrR
82k3iVJsVRpQ8x7HUZGUp5hrV8vi7kBa2yZd8e67BNWR/vCNWAsgbbqx1MuZ7MK/4xJDTgPVv48q
qty4hcUQ+dfok43IUJmcDNNhHoLoKSWGh7qBq/STqerzvRsgqZdoGhnmJlX/owfUnxhAWZJ/7g6o
lc9Zy5DGca5jyfsN62J189/Yy+NIl5kjWRLiXy8tImu94w2I/wSFAULhOEabuzPmFRTyCQu6oZj4
3jGn4S7NGNuvo0Z12IXivpVtJwEc2jy50Omclodfoi+9KjFDsLyiuFcrmd24x3KR3ml1duw/nZAT
3YMR5lDOfOtCpUdENODBSAbLCmU7u0KU9Dm1FNfLsInBjCU6keg5DM+lpClBMnwpQXb+sHsEhm0k
vGY1LsyaIv8zgDVMh46w1ZXQDWJGAB472SuLmBTnsYkmGJ20rDqF+OXztDfUBybaK85fZsmMosAK
Px0mcj4qdrpJ/dcdY42mLdO7sjRrsiwZTDZk/hhJ4ibC3ws38BysSsvIxeHsyAMjkgwFix8k8wkI
UdSfrNECcljZLPHfnRJuDAZ8qhLOTKkNsRB9rMj/0UfXjjXsd6p8+rvkRbhbqgUBfDiMwWxjZWcr
WC1rM7V2bZ/yhE9YHXXGydZIf5HYt2Svg3UMXwtf8+Q6vegMwXC38tYg0lsxq8c7Xo38mTaBtCSu
0fOouKonUYmN2NCMg0z2Di5Y2jb9wwttrQlYqL+9k9G18qEMteGrpQqcdxJpsmVadL3ar+EHArHt
6scw84TaRDeEfHHhAgyPKqZ0oAbZEkwTSDcgAwAikEnkY3SiN0ICvYG3s9iXrhLw8JKMDB4p/9QZ
z/eQZFLk3XlPraprb7mUOKNtyWgUByGQkgWAGKK4hDuRGGIHpzWRuOqAfaeUQch+nivwzCsjf5an
OsJCBzTKCfcUmPUdLu9v9JS5307MMZjrppgfPGOvV18heMAYL1clreWAH8CTMc4NvxaF/kXBLt7P
O7Dv47FdfMJr9g2ifYDYP6HJrELRNvRIqBLVEuEOyd65JoK801Ql0fdHuekjUvyro1c34jqNnAgD
0q1qdfWlmrzHKfngABW/lYhAwNJp6S1tKn0RSlkZtZXKK7411JX+mk69/dzvwGzZ9EikREAU139y
Qn2h4Kx5HF2KGsCmenxW13o7ewv6Ix9xDV8QknY/tkSAljCuvZbR0ucvDWBGw0XUm1omR7JbTcrv
SUngbg7eewfwOU/K0rhVRRggwo2fB5HPkdeAWvGR303cylY7AdjilQuaiQIXs9owDf6vMMIXji6Q
HOTVSdhXdDWrI50cWzvrBcoyPF5q5c1nch13cdeRSvS5SHpckVFkxT5bxe9zLZriND9WmQ/Q1Q0Q
fKGL1gmzTLw9d1gGrNoQIlYjpPNsDNPy5RZS8emwQcb0Gu+UCEnsId6/Jen3OfWVG/n5gcka9Yzj
DRv6HS3EwSwF5ejGN1zWZCfp2+Caos5JJRr/nWq+Tacy/SLMMJexgjbDY8WmN/1EP5mzZaLEm0bZ
fkPrXnPWA+oUP75khHqUcVqRGV3UWv801qwF2cIKeJ9kDgsw9imQTqtYU3TjEx1YqGd9h5XY8HmF
bk9MK1EisokN7TZKg05A0hjj3UtJfQaqqVOA2kAm8bXXQmqTsFTF+Ccn9D4WA/QKXYh8UrBaw+lw
XstY6qNExKyFzT0q9wRfTS5LnjNR/+ypu67tUFEn7PuFToB517zbCgcD9hZgDXDN540JobDoEep8
zfUMvsJPxkTGUUXuRXvV6/Ziu3AN1cPw3yXohSvrl8kfWnGK+Ss4oVySR7YzHrcTk9ThJtr9KDqc
RvIM3rVRm62eSoPMwC6eNLELm+e3eYItrb4CVYjb2QRk5zVdxc5Bdf2VL5UNqmbaEYHf4bS7DQnj
eBk/bsC2bg/oBIKRhHTMEx0sej2Sy9/RYEaQikf4Pa20PDyMedlGUji7wzAlAoWkgA8/meOJGDLY
yBEmxD15cxXQmas2NeFw1UAoHrLpl2Q659iZdvVsVXAGGLpUlnItlebcuPeA5JgVCjCpkHd7POGS
nNAm3ViZkQB94cvPPFfkr8l0zqrcOBjPcpvA1r8OKpi/3cX7YxQNlKHk1opILisudT0WbNIjGefc
Y1zuF3lB4uldCHHL/ccVU/4k4hATGEgkgIQM3D/shjxzVEtnlYl/noywG10bPDk25j3ZZXXodcKB
FQLdLa7v8tYS7vArurnxGZhANQL6vKW39BRsUsvMKOXGpIilzQ/7AQuGMaaJOld5gqqmF0MEQVHc
jKq91C/L1NzPNDYWF1yEFDl1kcRCv3SsitW4EV9m23zmmk0hatEHOog6Z+UulVr0o9C9ZId3nPzR
XEMUkhjnNcFcBe7zH133nULrl8JJfLB+CPv27y2MSWtSZUekkUvMyCQrz+z+nxba29JXfoT7hGo3
3Q/Yh6PEQ4CSPFkoU829elERD1blyyp/NroeuMMqCEmdVGm2Ib+1N1QA4O/PGJwYPvQW8xAkAOG1
zj1S61BsyICVwAr8HKuXELY5aSWIpIL9gGwt9LxZtmTmOzDhbpmTWcrHGKxhXmbSoXrgamMoskJn
gH1Zb+Ec067/9l2zTQfNOxiFCjasZ1/M1qV8QgEln4LQeIQPIFZj+K6YzTAyixnY0acn0e8PHSB1
v0Ahi20ViPH9V4apWdOanOfb67vyRQrMky4dqlOHDkAr8pnpCMegSZd989lPmt+ATKYO6yNmyvbj
ZuuKbmuJ6lzYR1hPq8RFHbaSVf+h3kdkj98+IZN+RieN8RqCr6MpgyklvMMcWJbeYMwMZ7h12nPU
3rzHJHHg0czXdrAZsak/C6c4Kl1T9AF1pnwJ8W/AzgVBAx8IpMEx8fVu1iMGTs7ijfVzGXVy/qYE
r0n0Wfh89d3W0qFJEFDLVD2Lba+4n9ebyXnrxqopvZ7Ed/Gotnwjhbc2lYleoM/OF/ehPL/d8riR
1Bg9SBF3P29/i7nbTdGkvrPah1WmIqMCMV1IF3TyuXCyzn7iPDb7c4lMZkhO+j9QEDiy1Lfv12cz
lZ9J0QQC/hEbHojrtycwyFi4HpV7T3AX5+6nsGo1PGuhwgf0W30CV5kmK5KODHHqwA/Uvzh0YoFY
vw58gDaBk/DgVji3shnItfMvraE8GAvNbNWe+ajaMZDcK/q+dvmBumcLHq/ya33BSlJDM6Vx/XhG
7jCsBDHiFq12ENwh8O6O0quYovX2Uwsc+knm2GBjUgTHRF8O5esNctDTkg3YXw6BC80E21beHmpF
E1rGW8SKVEjEPESkyeBcwHGbxY98E6e49OS8otKJ1zHLd49kzaQw4WySIOnpWNlcE9hHoWnoaZGp
vZLfKojiCbhmkM+TCaj1N78+3FCciR1Gqrw/HieCfeJc/RLKytAfY70wN9hb8SeK5M09TSNzOL5a
4dzE5YRC7O0elE1A6ZjWtMuxf9CTJIPAmSSVVmkACYsC8Q5eCGzajssinIBB1gkblf1n7jw1RRjQ
7US5Oe9M1qikQ/f1QfR4Nk1rrPPIFzcoiA2ozA+wzPq8XVYkAj6bchHdCdhitS+PejrqtFIUwLw6
96DAibAdGrSeJeulqPBElzeVpPbGx2n8BaJLnHcCUITqmRI4SOMKHXYNVl7S5YhEZdou2QQCmcyH
UBE6fy/a1yXGjWuM+61e/CiEeaVPPj33AHJfHV8UMXgrzUsbLDjMuHhTGSkqHkK2yUPKXRAOarr0
QBI3P8uGs6JRW2DB2kWgTyzOrPfb9hkNivSLLAl57aggK6eizqQU5DLKZIfv8Y42d4YZAZPHXRJf
pi1m3Y1Vrit12qgiK2egeRLNMdUaLW1jEVPrH8k8A7EuCrhxI/whZOy7TPVDDTMFMlmD8vpAZ/RF
4mHuP9AZu0w1FPMqp96a3iJaZyDOf0lND3Lcjc74x5cY/NzsVrCk+jDMDwJ1G11QHsqQknxqupdF
viJhiYp4nBgtOF7F+V8YbSN5svwjXcLRuGT4YURHH2ZNayKeY/8XfxxXXjPf5DOuVfKkJRHRQ3/q
LIJmAk6skJ55rwN736v/Q3q7BRVadYCC0mOStsd3W8txA3mJzeWWZAp6lPNbsXIJC6SkDK3wP3Jz
t6kol8W/wmEbqpUdmGGiJNG39CswjK4PSMJcyrwGhn4HfMH+YSI90Li8n61vNLpfePsBwj21V23t
kfz4te0QvjuJMVZAE2HSUwC9RjZw92lh4z9QtefSPbkFIbzU+4ibGNv8lriaEqgAL8aaD96Qev7d
rt6UI5JuBkai+Ijpr6wwzGet1Y6oPKcRkF16fnDOJQbJeuNJe3hvFhw/2bqpDecFTBw6+GzJRZ41
WrT8pJI4wpZl87y1BY+FCNQYmEKXq5tavP5GHI4itPf5biLcL2HVjNHzVjrWltcDSj/AA89J3ON5
lDo8tz5JnghrjP1ruv8vzU9N38M73kHP4Db9U0ZdwaYiaKeIAIvYYI61qKsyCy+gmOVAiG2nFPGN
DL9buKZTAJxS20zrrofjdg5RqZkDyFh2WOb3QVAWwEzFEN8QmDupj2YHTRbGrKeSJrxJqCac1w7Q
122Y1NOH9G5EU68idMNOvPF5Dc3pl0m6hjtmOsqEszClztQIre9FewUAIIXgPah/mzTQXHwpkBQ1
of6IoSjqAiSka/UW3vaze3CqNloCgEsUbf6T4ha667MhjWPP63nRvcIldrvDuGtoIfHTFg57LA3Q
QUt0t8RYaPNkw7UFX0mcxB6GQGJEiNqGW7MV2+H35YAKOGe35LJZGjTZYSqYwhDTJNzxXjdrRF30
CHhErSu2y4o//9mWK1ehGwA664RW6zBdrvd2t6o9oXZVDuLZmgtMkElEET1NmLm/CQ1GzsM4yYWJ
nlRRqjviq11J9TUfEiHxHNvQAgB3Vpf63oFsDBaQx4TXAFP0z8hQwLLnQOXJVe4mKv1qCxJzzL1E
/DdiGjEoZ4P0AJiszphYTQ8aEyMea+o3l6qsyfMnZVByxOnXcfO02cHHgRIxMcyNe1FpYIn1ZXas
2IaKN9DzLtCUDxRBNF1LQgCeR91xYqRDLjboXWJSLdewkqtk5+qcWvpjEiwXvYHeLKRaBjqScHKm
bwcAE3+OwTl787MdJs1TSye7BtTY7LIkVUTnXVtnilOEu0R9WkjxbUwOHl76OT+f2MjYZuPIzF40
sCsg5r5XSpuAduZt+/t2snwsUchGp4C/Pdh0usxwtpqHEP0Us5MwSbCNsBbQFI3W8AJFqxLU8UJX
LWVraWe6u7IJrs6Pk4GRAmas5+6fBtx6eTjff1RKv6/+loqkmY0xFSl6A/pUZy3C27ifTrrUyqp8
CtPGkETDwi0BibdHOG5Uhwl8qyumheNHxGNLSaQ7SsRYzB01zuIDSFDQNGW3iMvTIY86C3eQBrDs
WJnCXgwv2tpyQouiigNLKF74yyj2GJWSQYfk1+uk5gTXfyvaB5oWMniMvdb0QjWgZots1R63vjgK
pPnWvQRIeknb8hQRtfMdyQqs3JCxpZTqcRXkeEBl6E+HvDrSGGkvZRNzJKABqvTlayoFFvQaa7aN
JTSg9dA1ocw5yKKLVFukuiFZXB0rDl73sAW2i828FpYPGAgO3FgtGhq47NOcXo/Nz5mesgdgitai
4yO2QG4L4kdrWhAwgsfXpD/Rxs4z95p99IOQYS8nixyEGm/zRJpaZgDu4nungHs2zPlOXIeNlfxc
/e5BIxmw6NcDPDTlsYq10T+5xopKD2gEO9fgQuhEgqcRMve5+rAI3p2M24WFgSvteONN+T8Smour
lChydQYGDBDSzxCKIdimeuM8ueH5wQCfzQTjQ4cYmO8GxZ6CKTPrV0sdYyOH6DNp/We5/Km0pSyA
OtLeEgW46K2G8WyglHC5xPPIqlZZXotckhlQLcFdOKhdavdA0vFM6Ud14ZV9ORj8wNSl76FZfvTu
VHVj7YMgpys+ipr1RxmcXjx80G6eg6U20QFRIVWg2pEQp7e/Q/vvhVHlWpm/K8cLEDjm5wT+h1F0
axLjSF4A8C7K8vCC50h9Gk/IU4TBgYcqc2O8nmZW7L4ZPrcnqkVCz0eAdj1kEjzLCwq1u0+O84XB
6XpxfSoqpKcCMZjCObRY3BI9A1Q+9qTvarMyjXWNGqZTIoJT+SKGKvpeRADKF6qluenico4TKOaN
t2M9a2ljuHtT6ckAIv9L1Xh64f3MuO3za8sKmyZ4iw2HKgurX8wy4ngm7pQuHdJ2iTq0SYduTzbI
pc/rACLX4o6R1QrVCrCXl5da6zGI7LF5+2r+e5WW97XiLq8CgaSRYTQN6JTr/IEie7I+9zKKFpCl
BxHiM3T07fzJ2ggMKztABmMSIfEc0GV3diVPdHbfZQsYFhgSfPwJ32B0BvyAGPmHYwn6lsSzi4tN
YyGZJ0fnrWF/4heRecWZNauBWjZz+woAqjCZOk7KJZ0cSaFDBydyXH3EPC94xL4K4QYE6lYGtKQr
61+Qiz++TEL6BUEj5/G0XmrAlrIDPpg6LsjahCoCMiC1CM+N+bTERN4Ty7FYm2IyrrfpCdorlL5Y
v16ItX26SwY12bfy+3vH0QAUoqH+NE3gzXae6fY0kHwGr2/xtYSMP4xrRAQOL4xmHCFC4L0lJD4W
qtm6PKDMXIc722w8uFzxxtgEIViuph4nbPIyXYivAx61jCUds1dbAWXMjCfgWMroGP8HoOEcMCbY
aM4W+cHOMuk1UuAJ+MgJ4fhOl9E9Lj6oDnakKS0j1O7QZDCB3Nanfm8AVSOTrULwoUF2dHqS0IsA
tknuVq3Grr2ylrBQKIqgcEEIg/UwZxryNjwAFs6Bp/K4wk60MdrS1xD5sk4VjQ6e7MilBrhCni6r
NlJYTAigMtGbChLW8bIjIugkszvGmiFuflz0vIJQYY9j0JB9pQD8GrFFmxYtF2Srqahf6j9IM8de
aEKjXUvvgU6HtHmgAgAMSicTOc9FiwQS+BH4tOm0Dwz4mu0SGo5PEJR5RQ1CR+ru2wmvAqdMv5Sv
qcdzzLUdZjeP3sGsDIGWZZmM+FB7mvvmuArURAlrj0fIn61cohUsmz23wCRjIklrURt9YgveOINO
PHM5FelOg7oXhzOvgl/0uI+bHcSa7/VY7I5fKVYHViXn1nxESfhzhuDdu4K19zc+Hwm5T5rkdYJU
bOJxKOJ1oJ7g+yUAFGCw4qXiwHFhbSeUKrOZLkntYAhvZxs2eS9UspZQHMzwcbTSXpVdoKi6BNwP
7YZhbt5pr1fa2kXghOvbiS9pGSJaF4sTeGfhMwYJJkGlaxpg6jBujd0hlyDyTwk30XfAPHrFuGrX
guehP2LOhiUj3eyFmoxLimJSl/JBePlLexjIpGdC/7FRo0GXw/Qn+bZseKRysxVdww6/dXTtHmvq
kKEAI2r/k1KaBvol+Ic6eECms0AFFR6Y3XbEeTNQ9dZ3u9MzBnH/zW6kRXqnRssX1ptgT66QSATF
zvCU3drGrYdQqdaFjgm+pG3bsJGli+nMWrcfdvxdQCbc26MuXYAeunodOvkmhU4izU1euH7zIiMQ
Ck8bSLlIrsWNQ2IEtyPLLZVbjP1UcYjuBtLJcwamCJPzleOwjJYHZG85D2Z+KOpLD3sE8nEHUVFp
sFXngfa7itxkUoCi80xqNNiY33GwUYP/PzAVDFWLTA31hNcJ0IGbeTy4LRGabCwnobFzgPs9Eof7
zkSsf0smP9oj5Z/RywF1QnSxRKm17wDPFnzlFlKBXB5/j3JoNFcCNoFv6bnC8HwwL9+AtVnDp4g1
7QCrbHh7pXMzqnem3n4HNQp1OihI6JJVxB4z6HphSMzNJzJqbPIaxseLGxIdm0ePfiftQxigqaPp
dQU+k+LnbseOa95tKlE3p8L4j3NYKw9KNEypOGBXIVl9tcuvh7i99Q0P4Ttq+/lhUEGD3qo7B10X
jQJHC8e7MvYa4A4GDnjdKQ5BKAOJQ9jihpOfm/gbZiyGGBGSTfpS6JdyGhIhoDWsogY8HFRkvbtj
lJc6yBWu75piju8UN3ik255XbbvPxGAYLlXiw7p0jn4NLePfCYVp2Moc0CjG+szeMHr9Rq+x+ufs
Ata4FGXD2IuAjO96XRE7C5Mqli378P93IdyUEFYxJG9o9jzljmd9X+CjkzJekZ8YL3pPLcMrg+F6
pj2YKLNE+baX8OgcGDke8c/QTaKAPoAW5n6pNeSuyh4miIFagnUos0aYP8uRFykK8Aifz5t14M/L
P9UsGWukt+VC6RTcShTcCilhTBPFro38930eeVJu4MjzPjGB+5bXjDOtMunw4BYLdSFn2tvbspMe
WplFIRxDjntEtZTL7pSRrnLe3Ab2HKjmHfRqbd9SvOtWATI5SGVBg0wuq0CAZJROWCjPzRNI5kr1
w1qaoiU2jy/mE7QPY7nImv4vyUvNk9/4Vy95+qxHh/0yiqwXi+h28hEyMKwDVh4hcBtu89v1e8vQ
+0P7uPSeRSq/OsL1+2KsFGE2d6P/yJIuHqw2RpSS7UKnZO5VRnRGHuXnnjwmKBzpTHxPRNNRrp2y
r7nNhcb+oAZI6N6zZ45GWoy9PvVXOcDDUvpS3XGjwKqz1oD8PRc4VFj2f/nSGF6BYqgFc50HwYna
5qHv2ZQA8wTJLw/pHJJB7xQMcKVa0PlSaqRFW4vd92asn7je5o2hl4UdX151eQrSYto4X7rIVOf9
yezJMcyWcO9wBvaxDAIAQHQcI3DJ+XxW4yM8oA5zpCF9vJKTlN/J0IMu8h23osyMFWuXmEZ7Fdlu
s7IR6qvoMoz99mU7iNlQeaFmauZf/km5yvQXoVu29djhej7zUCmPmD3i95vew7+IXJLzat94pdPI
49K+Tlu2P5oyjcCBzMQ+0FB1WZmt6clSB2YuqV/A6ueskvnGgxqX4+FFruuzNKzv7kDqAg2dwzDU
lL0cIfMWnt73ZV+tqKaSwnC55DFSjE56OsxJYqfymrL6ld4GcfSGmpYOra9r0vlVrs3j0utI5WTR
vOlAoOd0mZwegMhyXDvkCyB++O3u3bBdHNPPlnRyEhnK/BXHW3cjRElkRDjeCZZdggPUXGkw1RJO
pUNM8Ca1DepidBGjWN+icYlabPSOJVlbROJSdfkUVoaY3oJJxf8W3RJ/t+xPaFT00mbzLBzaechL
hFUQ1DiX8sP/c1SFWmu0SxYf+7nczH+ayCw0DHGjLvSAs3jAjP1JOP5EL2NOM4z/THy/C1GFPawu
ezVB9BpQ8Vq9qepwd4uUKfyd9Tp6k6fwCI5rEuvlmljHOfO/giLAvaO+gehEWoLwxBBCjOm1WK0E
ARSK9QGs104nEW6x7yWZQo8PJmSH9FZsLn0w1Ch3oGeD5x/nrqWQsKbMyH48pszY3O5/MtkgucAU
dBBrHsUCctBSLobq9tPubGBsO9gdpesB8jUjIEe0t+1+NBhymgdhZbAIQnHbLsybkFqx9NfFFM20
CuNXF1sdVaUYYKsbnIaikLBomslrOPvijhi5tbd7v2yHRBVK7mOOVoJqbTBmBaMI5HnBjzulnjiM
k5OdNZlJqrJpOrxXhwOIZOF30oYmqhZudJiir6+rLgyVP6fMHhYbFjI+jXioeRTXyJ+PlHqToKl5
ar3zeRQJl0jaBUdiqyDOWVLsX/SUT6dDw+HahrFWc25PsBWsgFaWgAzFzfNtub1jcy9eyRQOvz3f
0+W7FoiM0yJmMiNYbFXuUOUzTA2yOYZpDIK7dIcmhdzfJ4SqB3+cGEqppyHHDOjUdkNtdpTVHPel
+A5LH8ymPMl5FwJ7PysqvYvH+H9hY9B9r1QE2VK/vpaA3VfK1IRbNW+A8sXuwrekvv/zudBet37J
vsp0bbg/nC6xy97zlFwMlLm45bLG9wmXZqOaAPcMDR++Vd7xeR3/mcV1f+iMimbwO0jpt5w7zBuF
rAK4f91ZiXqEO1hCROEjqC017CZUWvOE0NDXqZdmS68dBTB2ee1u8zOl4TNEcQW48HeKdRK0H94W
zGQnaKXBXpSx9hIk0Zrph6pZmuMo0pzt41Y/NuZklespKMeLmRwJVAU1YVJBkKC4nu2C7WjfTDXI
RMuzyARTAhoFo81qRSafHHbLY1V2fzWpp6dYwM4MmdhTUZIHhdzhbGcKnXujBCySm2BD5ZW7ZEXv
4JVY81n7PrpONI/RYvceGDJ57MP9j6PzRNqDX7e/WIvCcU52R92Oi8Kl6KIg1vOt4Rs5ZP5DiT5a
FhcS18O0tKy+gPHDyciZD9hmgsxcFLNVn0idcPow65erKY5N/Ld1Esqc40tj2MmtMBoN0UsOAgj1
It/Y7+8TqIZ+JWz3XGoiUw1tRHACOQ9/gYDY7g/TuETntLO0HfMWML/y/jsJa5AElVVZVXDZC1fi
IHvH54za7/84WrxL2xWz3klpWaYK9IMamk+/TST3Y73v+NNmqMCCVqPXNrrNf9nS9EEbwTWiopLe
P30dZDVX1sCqLfWhQU5z2j2/DLJM5vatUQtWF1fVAKQ4fvRmjDXFSWRXcdduWYwWG1X0BIdSzcjo
uPBAAK9w/xjgVilhY5wNtZy+UlxZSJenLQ3mqtYzdLUgVAn9tdbW+leRKLJSO7gfj3XrUfTaDKwj
8Q8L9w9ktvhD+jj18Jgxen7t47qiQmXGJUJ6HnaCAZm9vCPMVnCC8HqLU0a54Av22g7Ph96GlO7M
fyJgoiKm13xTi4jva3NcHeWzyilGxPU/XWSWzNG9W7oxhfVQxRy85h2+2ga2YZ3k+mdbixhQyWT+
/JlKKfmvDOESjrP4GTdnT2nO8ZZwmQTGNFoMKXQsuH1zf9DI1Z52YCuOMamFtGGZZonil9QTU3Sg
3NHaZ7M5bJcTo2eCw/yUoVfeZqs6DQlHFlrpKDDQB/jYfSCMSwYC6LsofiydTquEdi2f6KC1qn7v
vx5KdSOSHMUUC0VMeNOxxW6Ehl/ojNTkg2SPIFs7FQ6dm4pOGmvLIJ+BwhNvV1qYdP5n24HmbJ46
SKlDqc7SKxmTpPehQdX742CwZf4WRV7+2FkmoVriJ9r/paoKJm+J+pLI7OorMXfFjYSnwyjKlnr3
0PlBx8993QXAdMGwp2opUH/+f0apaGS5TBdoxdbYoRdCyGrulwHt0Xu5GJZqjg+iH+h9IXuPCH/q
vBSIFngyVZH8SGJvWCOfGjGUv9DUd7rTNsBfJfVgaLGfF8WieRbNolAQTOUSifXIoeM2FHoIIfra
N+w3rLKluY4qCL7OkxIDdVXbhYgevGY2GbgQXfKMptCZucUFSAnikd1BMgzQ94iICq6C2sIkhhfs
TIFnOeahPxkk1sT9/Hwan8klWRjBimdg3+JDLNoCYgOdgvmwVa7n81FjDP5G3yfahOdZRbVk3Os3
X1xI4YfGRkO/n92Iy1yF9zpbVvv1g2iPxEM7wBK5bTsDtzLDZSPnS8+QXxmYj+DB7ZwAOFvTaztB
hMOTtcxR0E2oBFjkTCuOuY1PAVO7jUq+Aq6sQgojtLzvCmO1vfiONrR2uFjAesbH9ShzzAlc42qI
/HNAl7wnUpyCiqa8p1VERQw1G55XMS4D3koe+z8C0vDh6h3hUtorUzPQOJy8B8JufuoSG0JJICvR
OBS796BdiI4RStuYALOy4SVSPAPRvtGVOwsnvmoKlyA3fGqn8UYcTPfP4m0bnXUZE/O5BcQp5heM
YVIxJL7XshjdUJ2f5f+6E4B6rSVKT3s7eS8eMVNSWdPWOqctp32HrwjSbKWKO88PLw6O7C8diK7W
AXkbcFwHzqxnfzUa4UbhgwfqUN+W8D5x+1YLEDZsjUbqLYtr8K3+B47SfcnOoIZne1ctDLI4g9oL
l6WAu+EaWbHurwdwPpdnp2IlUYKwdKCS57o26nu1v1M69tHj88u9DzB/ceeSGaoOE/kh827jxYRk
/ktWfXef2QTaOU3wZrFDtNt5I5x3WHE2hRc+qbr3nLCaxMv81On0MzK3vIB3Z63AOWhLjBtattNn
iwDdJClyoganjiL56eh/Kan297VjZIu0Fi8o7JkPp/z99Lipa+GytwJJ06LPoWpAFX3IKqj/AX4q
h6PLDAugz+BFnfzQ4stgyIogrZPrbpb4C3350wj5CWbWzGfAgi5vpfPPnrAHeVHMimFXKmnU4QIG
RTIc3bMIZAOdS1mpFs7fMamLSpy6fFadyJ4ixjrPECPpXEuwSHFa225vmiYADkX6s5pJdgGIPz+t
G3MuHAXu0wx3Ug0IiJlruLjlqUu/6a6uBBT69pNOB/zTfmC/OgNhyv5D6iqTTAlHfwnWtqTANk0o
rJmTxQUVO9Avya6kObyiTLGgyq0VHGymyHFetYhOpYdYKNvfpRlutzXbJdUDa/QBU/vHTkBzzV7j
j7FNSbLDtLRMKohMdtBj9o9nTmH5nqEnvNWJxd7zLJPdOhNOr01TCKJXQB4ziUa5jA8nOWqPvR4Q
RynUk3iATk2Z7FYQUlwupxp0Xvnf9hip5B5Dyig5SSRnS75cZFV+LMKN9/V6/v4yvBNMDurVy1YF
pQop7a31K6oNrt5RosXtp4h2ljBpc7ywa64a2pyamlUEqWxplDYQeqcj0sSZ8MichX5gBzK0+deB
JKJ6b/6SPsFHSoWBLWsXuZDOasy0hob0KuiPQfHwKu6X0LJD5184m5RB4sAqNVf2bMOsNESbzzwb
1gzD5HwA+P90A7qIR3dtni6OeXAnvkTTtkydkds5hEUEw2IV0bbvsdm3UJjZw+WOiVBKFRdy09HB
VB/fET3vWOp1PQVPcUdpIHZg/zrMF2Q8Lk+KMVp91M71/0UscKh3MPxVv+pV9o7C6DT7+AbroDsA
p3ehJiOZtS2hmYjUIRtiLppejTelWZZmOTwMpE8zmexNIaWpR/SPDTzj/S87SH5qEoKk8GrKT66P
IRxSbaGawwmUngnL6nQcO9ZZ1heSXAn1vvnCF6shOcMRzVJnnYZwh12sTPlXXGY5g0NaFFSqSzrb
lId3AxJ0Uzshv2zd7b9nEeLym/VugcMLOdN78gI8lMOeIY6vdNyppjiOsYJySeNpSbiytl9jHAQy
T9EXzuCRkwh78Gx7UbCG7DnGiN4U8k0Rz0te68xElpblYLhte9I7noawJVXeGdOLKGJwlwPI7NLi
4MFGlVBndhpTkymoJHe7NBQuYr73TFyQXzNa6DVg//K4Z/yDNGqML4sdax0DlSCry28TQdXkbeOR
mJGlTATPuigVqafm4eoI21N5zBBiqLD7JiFWJQmDlU/ocUpEYrbTvc+O62sw6TsI9+kciKHR7qaW
eJ2lSmXQZSQqUfaPyd1Bd7rG7/qWNjbGkN3kiNS1Xg7vTi2O1EHUSfhy0W/Eygt8dI8FY1tATY+f
PbRg1jJ3jfXI+4DYYbV3+axa7gUtIApUi8uzBbxqxvoRhWZzTLbMNDdI2JJxhlTFBoCR2akgQwTn
dEws+81Wpw4jaQeOwQuikfT3q8fvark20iSXW30/dvnF9mCuot7q2EmODxhCxnBKcZ+zQ+48cXCE
ne9zFaSaFRA1WnNN6oNWoevRl0g78NKFwGIDr7EMmZOQUpNku3V2YIrx4dguajRZD3MDGAejN93+
+5lWccZFkPOaqGLiNPRAFYAy2031A2msww04esOhH0HGZVcQ0qNv+aB+13awi7R9reijFpqTQRN5
yutPFxS+WcKZJKfXs+TOkpVWWvWsx2UB1Og+mK9lN+fpzMWm5FOhN+lG97Qe4uznGHYZCjlCmDvN
fDpYDLJnHaiBf/f7jnWwviGDDXwkYk9zLmp+R4XEl+5UWDA1ybZxfsAJ6h0GOit/NXIQUMjMMomY
7FEBgPJDBQv68ZZmk66e19tiKDkqPHp1AW9oTIxo4gcXn5waogzfRgT5ZvIklKIGvQdcVgLWYli6
Fwrnowg9sMnl7YSMhMalWo9e7EVcA7isQUWgdfE3fVw4A6iGVJCW92Shvki/Gz5QChIoeP+mSP3K
net97QrPZgvNEJRJwqeqm9uODi8x0HhTUKoEs0qS4KDffLIR0np2igfM6Rhsg3u0dLuTzoCSc/rO
yms6lde+lkEp8JTBM6Lj5u7oVGvCwlSgWbmv/fJKIcJz3GC+AVS8aqLo1Au3FW7zqIFqKzhlLt6r
H8IpDcF19FYcQu8GUlcINlxWJ7TQnjhz/R57NJ0SH/OTJT5GCkpnILK3To9uaKxdQ8IAx3YloPGR
hu8Yq09TrtzDT7LsADyP8nir22GqUTrFrN8YcgA/bWPGVmGmwbrXATjKGeCt7MTo6Du4+kJhhKSF
MtMhMYjQuNyjRGeqDKKa3dmdG05MuTKZoWrZ+UGjTqEIonsy0nBG9m+VzD01Is1sPVbOmuhLyE1c
UTQjkoRgTPP8avDYix3kiPiTXnfMLFQ3DJ9bhByFdAjKWOxzKszjbUC0Vufdt23H+Wt9RZZrFFi8
n5mJtphFoEc0t5j5q6LHTaW3ruCqesK6Mh8suCYjF/TAR/a/ZtkUQS/7I0R8UMZGx58euK45SQG3
DNYhCb6UrDQX43yqNv/leuih2aohwxDpvBD1dw4md41AE7ztwH9tiylWT5K8S7M9X/5GROhtTa6V
BhUmEPG3ygAX663+dOcDHWW0TagOpEArKRSfhuSgeReI0U1NQVlECi7nGQDT/zq46NdyMSut3Q3A
QKAURMKH8I5Kv+U1ALgBU4/SyBM/Z4lDFwCCGEriHFpEetiMek4jAIltNaVokYoh33xgZkONnKcl
57KsF0nQhBbfmtwUlTFC5pTf2fTQM+H1KD2RAxEPIDbZcJjpEutOQMZEIxPl96k6wGlbCpqppjD+
VOpBq8wl871MkCY/EDjvscunVIj7eFQLGparJ6PvU+vcqijXkf5B6mLq89M8QexviaRdKmK3KpiR
bkqVGFLFKI7GQ9RLsKHeVa7qejVtgWDKs9iHXKxoLWkgzhG7dIBY/NieU4NPRhrSEwYQ328E/PGw
PID2sJbM9dfLVwNiu4BGreyWNpfdCPN9wgWsFd2T8ZE3Z2j2GkyqKHc+tYW0uIOUMjNZ0J/l9h0F
gipjWGBL1ioFCeTcS3Au1CodeLoSaOMHJ+9P036QtIjfuYDxo7eVJqgVXP0o2KB/pCs6yN88HjDF
AHQe9n6ws5mxERQGz/30rJxRiHgbmyTsd4QU3L3cst7uE6OWFsnyP7HUsl+Jql01RCvt9FF9o2kk
EKeizP47ZQuIeqp16WIFyQWLSAI/rFVM1Ue9xpBv8/WHcv0vlsri1b2W+f4+VuNzkw8O2MvZ+2TQ
2OgNDrq0zMq60HcwT4zSRz/+M68nC+/FU/2OyLHPWRIO98J+w3P3g+ycALL1qaI7SvosZv3mBBM1
bR8+ZozQq8lKbYWpvpe6T+iWsaI7pdWr0Jia8tAFX9V16hyMJOJxBIzHv3WO4/1X2zskTtnOe9oA
iSrmzxwbNwGdAVv7hfE14O887nm8W21OkHVYui82SHixyJ3ck9Nx1RjBT9kD/rUVMzH95x3BzyzM
Jxbi5BW1LmuxiTQl+5GS82EGQtqt9gYcApfJ26YBkGDbsMaa0TbW39uctQCPfDDVKOsUDHQ05afS
JOljOAq4pSiw6Eu7LuevuCFxW3qr4TABimpZA3KstmwZg5Um0Yjs/+p4Lr+nFhtl/SxzXDT1EzGk
mvZsuURMqT6PrWh7BlI+5uUaWFysYDhHGqPgJuwCOFtRvODuqFigYq3HIw+6Vaot8AzTDkDZJZFw
zBfmi402r6kxYulgidwZM2MJSBqZIHLUGNlxJdK7a8CrY34PWnPC3AuhqJsNr56B6KGij9D4inDp
5anaCrS/YZCx2CSUGJJDKpTDhgAwksXx+QFpi8rvvBchRXCMY8esVFMj4c8AMEnoN5PwmAI6VQm/
rEwz1RKbg5Kz0l5QueHXo55l0oRP7a8rxvqD3ttz28Eu8sYfoQSCRAMnn7AMzFnNrbffsDl4kTaa
hGTk/tkweyJr6GT89Wi06TsmnFfw8Zb0yEzn0szaJGGhxpFRE10jT3eCejjZOLlmVi1ZF/ZGxoCA
6OuXveauIr1zEWjvi0VakwecTaQFf0a9NC9fvIS9oejHCP4uJJ3xffV0J4DtDRaQcz+bl4UzOKQ/
QEYDTrYJyk0VUS6RZoTq8Ahk9vuxhpHL4bR8gINny/6idLccQDxEHsP8EQpF+VyU3MBW1rRfEz4j
5cdKZMtB9RanWfrq2oQVZfkGKeYGMJyplSasZrEw/2xVH95NY83TxSF6CblAI3rA6OrouSpQHDms
ZR3XF2sYAs3Jrtr3J0rpl9KJmKzVv7Fai20yzNAQdQ5edNyT6qZGq+A3/lL3DV81S5ZGW3aW9s1l
59PbOwSIHaJ7cGD6T8zm5v/axmHdSZatv6aVWLW98YqPD7GWkB0prbNgnb9gpLnwdSmda/wpFWgX
bkEgFWNEJQPbRkDVWicXuNOhJAvjEyoEJ3r3i421r1lA1wuqnk4AVhrAWoUlf2dHgc0bCeK3v1R9
Jf4ctKZAocbpmi4GuLeRIbYB9eWtKeyuoeqtOjxy5CtGH4NKaGTkUsbPF0wkhY/goSlWK0sj5Omk
ipGCi6m7KctHv6TFUiAMkYZp7fVjgq2kATuKQ82wAYKJx5aZ2kYkxz888O1dyBkTtw/v2pmSZUm5
NoilKCg9S0VaR1XURJliA5h1wBES6d5WCXXEYaV10J05RKQ8q28t9qywPtxP6/VLorvJEpdgyih5
Vxzdp/+i+pTavnwa1GNiJZU05BvOxcB4G+gdrhcCjKqIYMo8jQxsZ7LG9szf25AZfNb4oVZ+/SEf
wECTNq4eaOPWiAollDRvKnlrsg6bfuXFL3b4kTIjkscEFUhPYMeGqvh5HfYqS3yxgF3UBvAJWF41
KggLhMUeHSYw/7dKEvUWr5LiIsP0D0acHp9AM+Ih42qyZsc+Atwozks1pgMZ14I2fUE+R7d6V/07
2riOIXqH1SOVh9g/XWnelLj1Gd8wgfqQTHjH7dKeaLrJnF4wMaO9vG2SRzNjXVlbWOGmke7bxa/O
Hk0Y6RgleFyGqa+yHTSpHMaEilZoTca2MNU3BNMGqSBUFZWc/KgwGHTDqN36TSflNmL7tyLARy0i
F1Aq7wSZADh0nYv8ARr8nQ3DUQh65SeKWf0gymEqd7iKuthLHhIFfJ++dqL7QaCTutaWULXPKOQV
XJrLwSew7MbruC5fRuIprxgRXKSLnwqmDT+mCpar+LcAqGIlhqnzYmVKnUO6OCxP0VvVz2li3jl4
CT+JjLIGw+Lg1WGGGzXDv+l6cqZ9QmKsFUcBzrpBE5zf8gVJIrIfsquGbO4pnaNA2GppVziSFYLw
52oXURMqUsJm9ePku/lmPti9FR5UdCFeUfPecCYvJyblzJL1t7ERqOK1jOCuo7oLNs4IP8Mz55T+
CCXq5PSWltHHHcyjNXOLFu4CXeDc2CnyBJqUQhF+GTm8TKhHZYvSfcdEMRJd1gcRuoFlnYctLf9V
AXxkAwFiTdplxWejExgpFY693VSEav7QxbQfC4Z2A72+w/nlpucjGlhhP77F8N/f+yG+5Y5wWV1x
FrLlvDE+WfdPaLhFVNUbxlZzi5ngng47KFW6/mpz6ktFGjVFAsmhKivT6cQ/JbgFfmJ1t04FK7h4
d/2aXxE5et20Pv+u2cOnB354sa2CHk2Ofhq7zoLozpWpwkIRsoVOLygAQd+3RCKWdTL40MKCWmGq
upZpBeDAKLVx/TSsIxaE3NMr3/D49l0ujCihfpyGS66yiIDzQlzx64kNE7AwCr6dagzUhw1LNxuX
Q5BZQxf35YbPmhlSEV+zKewhf7kdrEUknxOGWxyvue5Tof2R3yjpkb6sKvfCuZHo8+rZGSIjo+sn
cTGjLTyA3UjMQGjEo6yAx9Z6Ycqd7UYFm99Fj39aT3AWmYjP/YHEvQAm1RxXYaC+B5YfOrsod5EK
WIdrLyw3VrqF/MceTZ6sOk1QwCeLsXkrFGAiqklc2HJSiOSehBiLtBpE3jttIyIoONgE41q7/bkf
ZIhAoUwpuisKlnw/Y6cODm8X0cmW0gauhVh8ViU0ZQWsDzI4rG60bzxrdzT5vbpt60lePpHg5L4a
Yakh376+BU2tY5/hro8iJC84YU88KJ89uNvn3Ql10e0cfnM4h8wxgHR/9FGiLqy44F3+HUmnr6kI
2fYYa9oBOomhraulAjdxJS6wgAYtHXiCUU3roJxlo6dzKxOLDIkyjzjmuOjlN2EvsQltMBTgLLYO
K7xbuFdN7HX1BE/aK7Dl3zXbhqaicPq8ICgbbNJbla9QhCY2sssHKEeGymALxOdqJWSjtJf7pIZ6
1/l5SLtfSkT4xPH5Jkcq3EHwzysQ9W/1rZvf/SqEqgqkMBMD0HmZa5qxoqhZTmBnS+ShoY0I3RFQ
6LqPG8ZIrn7tmSfpwHBrojPX0MzCpl6dhUzpONo6daonv4YEL8UdytusllM88HnTw55nDQI4ZIaD
jrQekmwqN2MdLcVFfzm3+j17dP8/cKCg26XTR/Pun+ugd3FmataHFVSimIbY9qV0P6Z0GxQn0JBf
c7+HB4q6Rb/eQaeRf9TD3FNfDPtTLMvkMABOWU6spnSi8m+L3OV1L/ZsPM5udekT1urxE/gbEhU6
tILGMV197w+1xJg43aVG4Ry3vPEd0/T7FEBY+mXV7PK/DRuhq4TX8UXQIwJE5++4g8VQmHhor5f4
vpQgDels+xSbCsVV3eIqnyu3IJXen4xWHJniEpXUakIEokexKYh6ZvG8tC6+YCgpWaxJvsFtwhKp
lYooT5RIjieY5IdFw58tUJiQpQMszbd6WUMAicJqW+1JcN0Jax9n8uHpdY1u9+spnW/V6VbY6Qce
Q1tW+qluM8rry6a7OD1lHjE/GC4N+VaCLUCpnp1GF76j8KCFD7zCCxUMKCXj7/Nwht/+X4PSIvgl
fEWX8NUxLB+fQ+EwKRY7F1wuWbPQGC26f/kNH74cljwOboWP+WL/2F9NeWJDBJwRosvuifhn53Nm
G3XsDnHwUHNsRths/GWuVLDZnYN+YIXtjasx7gN4ykAAJAzKVQ/oxqcJbVziU7KGH8pnbp5PFwCg
nsprj4q0dzcsPdd1M8eALfksiXaBQemp85L9nRamL4lDfcJ0Dl8IfwWCW+PEZZ6EnG8toH7SCw8R
/Y+uoIC8mVBb9LB1IgbMVppsesBXY+P12o5Dww6xhmlSNon+Pnlgr5Xdn5vFrhC/lkkK4kUTKLQZ
831YMNlC84/F+JS3NpLilOcMpUopKA9zRNKqiaIAisCj5P1egxTDVVpWFPNXnV0oe0ssfA513Bid
bmRj2MN9AJO2ob7t2ZiOLlTdMsi5xd+Ge/y2SLAIrU55SkQoOE6bf284U2+wv794T/zoEl9ar0ru
agqRfMA1oaUAjK8vZrFmbicF1NG5ott8qQSO7oqtg4DU9N5f6KawikOkHcVsvc4mft4DiKMkYDIi
ZprCiB6AqNRlQ9uU5s7aACCdlwHD5MFXknqg4/AvRvC91LExIH2jZ4uJlR+N6zquevPsVDStJRv/
6mtKnqe0BWwIuzTogLFolbQS7P/OEXzwBHdh5Gpif6b6lXgYIbXutfdimmqBmHnREAAQvOcMI4yv
r+u5cG09UwfW8SNYoJFBZ/ylm+SXSSPFSbLa1rirVs3L6G+rG/m3oafbkiMbXsNcl/vRVOLw0t0p
lf/Plz4jJs1tO8z865X96P/VgNojWXhRUiC05UichMUn/8g5ih8uvkd3FGINzTAncrmG/9xnXHw9
aHswt2MWWARfS+CCVs6UFipjPlP1RBH5GFeU5Qr4RMioErji+Q6Tu+oTMFksv0lGSyXMjSeI7GFl
UOpXws2X+J8JN52F8ljr81z8/kZ7UYHxWDI3XsPdkOYjXmEpZFqgnmJIktkrn5NacFQ6Un5wIpF4
M7BvdnX2+P1BuxTsZ1UFb4kbsBxtyzfjuuDY5dqjx7NxaUv5xdNXMvGEiS920qDpMU0po0cu9//O
el/fh4cbGaa6a1qzGwn/ezuwhx0zk9PR+5Dw3s0TKVeOVVrGzqvLeXn4I6paK0TVbr7vaAPU6/ev
X4wdB8x/SqJIJqq6ovssKuQNpkNd7Mv2/HY8ZxAcBIa6LHou/IpaPnrwHYevZgf91McD0relKnCx
UY+MY7sARwGr0ltGKzvh+bt3PSk/AWEchO/dlPZLJi9ON8oDLdPYml+H8z2mxnE+4jH+nbcqWf7w
XFwsVm5xKDvp2xJZnswz8K1MRthQUnnkLfoBpwC/UQQGdwo+grmPsOZ1hIL8DbNeH6S6Sb7fy0+7
7PVrHqNvHoIwpFjCm+N1CdLzYPRbIU6yF6xBa7fASEudmC+pka2qR04gAHQnxJYJdeeTlFmQMzh7
+wt2S0jLShGGIbBOMVBFaWfxsHKR86GUyzx6+GHeZshn+pjgsrDofihxdLynS3hmZuWsEOExz/Xh
+yEtlPs+nn2Ljb5z5FzQwm1agZU1DIa0ZTOyVnMehJyLJHwaiCRbIR9MMPxwpAW40dI43Y3ZCM9A
i0Ng6BmaT5UN7daYwEP2fHl6LEkYaQyovPbx0mjUZxR/S+RWU9vvaL6FPLzuHmYiNuB+J3OUanvW
vArbLJgb1xgeruCz9sk8bRMLC6AWamLY2tcVwxSbUl0MWie80F8ZnrhP5pQa6RNIj3B3ONVVpsVP
6Wn0DNYaGmmSPIOQQBO56ilokx3jGXX8uZqwJkxJQC2rnwEyoXmC5OrPTj/p1SDFjE4FsnjbJJe9
Ixn05/6i89BiAKtXksGvoHpJ+tJe1a5QUyzD5l/eDXEf1IYK6hOoJB1g4nRvHRSS3N68O/qZXRqk
DGx9xRxWGCm7evfRV4hp1p7aujXd9GMGJczy3UBRrC3GxSQJgQJFNfaCNB/pvFFotbcVNet9zn3X
zsZC0WC48TnroGRiVRflhb5MLJc8MZYAEOTEPLipQiVJwVH5pdLXXuYppl0yWE9CJ2EsLhQm7Iiq
bstACF5ddqOuahBvAaVZYjrT3UBMMGM0m807AKv2cmw7sIPn+S410nboZgX/n3E5pRQ6Y3D/qA0y
srQZ7T/UCp/FJn5PMxmkpZfUySicwka+ZYvIsgdM+QOH9HA9JegOZFp7sYcrS/KyF7AM6gx9c0C+
Tfkaz5/X5Ds2QtfjjSuwWRR5thGlf8IxfvYU6ScIvCtHi9dBC6bbl9FcfhI537FZf72R6bVsIkF3
2GvqU49YNVLAiZYwnRKu/MaBfOtMk9YuuE0OmkKBQTm8DnK/R04zbJiFnHtRiH1KUproDBpDhfPS
E0D3DFnGLDC9V1oZUFANojdOOqYfQ+1ltvgoRxtFaeVkH6/wZQzMu5KYBkKIzKOYOxh2Bc2wEkTp
TPFaTvDMcct+pq8gVOhMuE/9W/hyrVaELvwcgvXfsFXE2gXE2plTJD4xWDGgHMQuAPxGL63zMhFG
0fKYJ0cZ54/ZSoF+xnCy9bhmyTZJDeB2b4Pco6pmVaeGTMbworllZy4lw2S9PXJcEg+5kSUB88ZY
LJbhvRKmkxbvyZzYAMymnoOVoXVQUXbNNNTAJie2mh64v1d47/aS5hj3SSXQ2J1LvW42J4DieZSu
9kS3AWZCDOBL6aUITrk4/iRNf2sUf+63XbtYHf2ah45SMSXKjTRCBHFxoPJCQGaNbPBJp/G85dNY
tmzMJph7u7DzUOABKXry2jjTM3iffBWtMpsF098JNKHBMkTl1TRdfSb4qFWSKFAHQsszEPASTX5C
TIsTsT6xoeOGt60qRMcLTFA9+Wg9BZuaGy8pAcDsjic5rl1YtAYib/qiVPpV8EoL02QU2I6gFT4L
OmjjpXU7Qi7i1JXz+rvA89/IkaEcK6dR+eZATq9CfEv/D0Asyko3hyF4HsOok0FHNtumnOaolX0I
fSzs7czBdVN1SqneoDPMtydxAjmh47Omee/3asz1a84lvePnTowcXl2R6iaPKUUnn01fvE9mbuaA
0YYRh7JXg793HAzxknN8APGdoVln1X/44COc3QbPtMeD1FlOQF3Xzhoeua2UFMSMdICLsJpu6vMy
1VQBNsBGo+a5Di8HeXuZzhA5l/gklSqRkx0oV3MJK03TGgoSnZOICiV95vjY21gltZey8k6Y4/52
ITDoInuH+wjbh1jA6n72lkrbUu5fVSKrmwdzQctkIFLVPVn0l67aHgRwVHSFfMRln1PxyyURgSQd
PG0ajdCU8JGEt43jM6f4N5l63HlbwkgqlM8z8R64WEh45UDHsYY0lmLLR0zVZuajH9AKkQroalmF
uusg74bGlkZypdlRx5WZBfHOaloSiwX49hE64bBVV0WXaZrdFhOdGyjinHolLZwxc7uqEOcDf/xa
iV/PrN9QrAvZy1rEESIkZQcYrNFz/+SxirgJ+O3SgtmHLE9LbmICh8G7MIBRBkNqJ9SYPOA5E2Eh
Pf0fbGHoFEdUEVQ2x3x/Yqj7ouLf3dBVwo3GfHPDahLxzXkWRn1pIkeo8IWwxn3jr/t13O9LGpy4
127vSqpw8NJm3j9wXHyys90GO7XZL/AikDzbuEoFnbvxiUoccYlnEDFHcSikTPKp5FbbkqMetROd
Ct09Zw2WfOVc1HYtP9BCUIDE+QEB1SUxszdtUeVUOq06aqNYKRFTwz5sNwgPq90H3Tyk9OE9Sulx
7u6BXAlkXmaN9iA5du2yxzbvdLZ8qgygeTTo/1kbOujBu2ibMScUhxYmJnWIQTtxRzrOtU5pTWm5
c9bEpPLVG4quS69PAtEM1d0sbsIs8lXeKP/tM/52Vyl0nKI/MwH221WUcOlOwRKUeDnk5n2BPsXE
F6KShx9ocdeFD1HgOWvqIZdiTZtr+i4OsIr/UzL90dc12H6RaPrnrFr4IlDxIAmM8RxbVvMzgxVQ
vX4FQx3DDZnugl5VZPGmJ5LvFap7V9pRh+KnJLpACFUSUayFdBgqpYzG9ml7zqUy58nJYuUSSLSx
pqxYnmqduCBKD0dqsUhJCfHZc6ciXW/DA910Cs3uLV6xHsE5H++C6RelvRzPwkqBWPsytfqhd1Tq
ZDQAj846iVxbG1qpy6WVSd24fn0HuW2xMWPxy5sr7HmSE/60XILdh89+ktJTpA0QeADNYUUfg+Pq
8Ctym5U82X+yfyV52Ur/WpYB2icMNYfFhJ3ibQFPQ/8msy3sTyrq8Kx852pORlfmN/YDozo0v+oE
it2634BH3MbBbfMh+wK0ubCEzZsSpjQbuSLjZ2zU4eB2q2C3H4K4e83GK6w40jhUVd1xuArx5I7m
zMzdnwnbsTRGDhs1EqTW+lZ0kpOfZyuh8ceVoKFifXhW4yLh1DaOkm3Tq/34KyjVfb8uwYrl4uve
XUA0aEI+fEeQKiMb2GakAmNjei2JJjOJcGdPnKYcEbhLzIiqTVojSWLY/eYZXMyDQb7iGpd4+Mdl
atay2NWMGUeka23VPzMPK8/5P120kx8htFZeFgU35sffL0BAZA7cVhCzb3TmkpDJEfCGEZ1Y9/TS
HK8NtDLyZZbz06nXh80J35/gZf9AHknb3YD2yheVSj0R4emh34dy5FKXBlM/PxAQX1JSg2VGEs95
tHvErXIARVmEXiAPIDHTD7GCPzmxh/eGe9YaMrlXnsKOmOdepweJ/CoLrWGCVz1ZGV2sjqCS+k65
4Cni7QBsE2JOW4qXwll4UJ3XHHPwUQVfIQnoynPBIo5At0qIQoYxomENktKNZT9/kJPXAxPDxSFi
2S6JTUoN9NijxFTZkNiMsodXtxB2r1Bdb+nRLQn4sCfwkrBJArNZjCgFDCjl4JDqhayt2O6B55cE
EwwJHUaqt6O16G8CPXcweG3ffGVfTgO23Tq4eDo60SNKMnDsYnlcPIKr9DR/zFWyt9kiWJHRtGio
Chr18gjkMQ0Fj75vqVb7ch87WiSxMQ+nvIuAmV/tiHljVszHmHXG9kjIFGdfPrAGn0HWDszox7h5
wNyXiY44qBOTk2O9EYUfqFRklNDJd025SHf6KHnSn3aQgGfSjkExG6YgtOlUnFShv4Zl589b9i55
Tjj7xnycVStXIlWBuf/mMj7e7YRywK+aObWHnCKcMLX+bv1Jb186G3APm/sSaIy6KIB7xSspPUId
EPbxM+ogQGEcuZaozPhy2ssL0DxBIYorOPx6CgPpZGlpNF1KMbmFLX4RuJ60r1nMtGXERHO6dmPA
BpYsC8gbInWomHPyk5RY6HZELPhJiEzawwLq5MseGw4MAL/GgRcIeVAIVDvtQEFcEuMqksdEh03M
Zts4w1KpLKvIC6a5Kj1Tti/inALenhmMFhMsQjjx8/MWK17AUsP6PZ7HKZKgHZ1flFtrhaVTJV0I
IKZQAeo6CAl8vjQVbEtyvahjlGm1rOI91WFd6J4ZPqB/e2Vvdbwr/ldigYImg7nqWiJ4ukr533mw
p9PupLfmj3rAceK26d3q7SmJ7RL0hMlwvls2Cg01ZXIIbQxM3irVxHoosh0XI11ryD+ig4oB7Suy
I8HQo1fr2L9LnFcfAn6FGux/Ow5Y/9joMyuPjILdSC+1HwZLMlXE2NPrFWH/xrL0KStPJ8td7LFC
TcM3I4AaSzkDOCgoO9fFOXA4bgvvbZcyby/Fdmnb2Eu75sGf1R0+aJk4Cco0J2IXvvrTnwgpqa5b
oZ11KuOyecikX3VILlfNyTm0EbAcws7WEF4N9IShIfJoTDXreERD8QjxRGT+XmSF3xm8HbqTvn9Y
Md8dS0tzORmTmwgAAQjnZB5Xj1p6Ku8VZEoHj0Czaa41QE/e1bpORgmIZXSpNNSc11NrXbQLfNgH
xCDeFOiGRXiixHLzK5/BlRAX7VTsXHhdYSntFhqAKaR3AaZviNSR2N2XFVcOITOfg1fvJHlUEntU
xEbkhpVtOLYoiF5fDqvLt17CkdOThpilEYSJFM8wRrtJMLgmS335UUPPV2hizyVEw+RsGH+Lkw4s
/2uRMROdfCuvNyJnL4PKeWJp2AnRIDeotaSRHgVNYG1hxUm+kiy+WtysidAkSyMOIiDuTYLrANAN
0kz3tDl8DsbfEezctWzpTG6OjoS4uE1MvxoR8ilE1avgkjlCFFshww8q2YwDag+zCvrtkaKb6Sdu
S8IW4pYFc2TDeG87+CmpvIL1CxFe0L3zawQKzfmVxUedtoJ4e90yOwkwkytx+cZu2aE7pCdpe/Iu
sWAwZ60QpMXJQhPuRAh1u7jJSGbPNAF6/98AVIApfiQbQ8CNQKZE8rKr0xLQgNdeh4lXutWe/o/c
P5teFASGm2fHoSKFd0Kx3tvCzOn6xlh/6TIZbCKblkmF8sV1I0nPMNjL7Qkd4SaQWxGySS11ngjb
ua9JpC7+XAieLIopSFXF3b0/XwCkt3+wyLS/C2G4IFrzodOEiawSt5RA8Xcc89H4P1b+WBSEc/EC
9XWoewtXTL28ZJmEbd6Pv8jorr9bdEFUYVUtEy0D6dDZwPz/OiHsKhPu8vQ1yL5TGacWDEDxNxZy
m6tY0RnuqsArlhZuu8GeKYlXklI+l0PDCb2lChDdQ6pD4pbgerIFBComn+KTZeaU/sp1mdTefh/H
5pjtKhz4uAjQchLazOd59AV8Y6siQCbnWDVFsfBZr/wSLl5uVA1rQKVjfEOCfEXdJtrteQRh4hTl
agGofTHLbUvDbyNNDXyEoVsOKVh5QWoly8p+f3Om3ytQCfF2zvNXaLEG6orjFkZhn+1GgWoZnUul
L7bW18gVrtB5okGTNZf2rerUczNTs3WBCHMDLQIDwiAf1xcE+Bfr/MErtvoFgjFLgrFyDCfBEcUG
qekqf0uMDmiT34DbLMxyuRfqwfL1xmDyJOrmgew7MhYx+jmE7sYuiCXYZAkFfzoSf6BgXNpSEshu
CVeRsGWWCpcKGR9okSmScC3A9a9OVGov8Iiw3NaM/MZWzsDd/yR46NFvPaibo5S977Zvcwf7rveH
+6uj5Lxvs+vOaAgmARGArrrH3yjOTVtoXr3vdYIrrtmoWct0k4BalSpI1W/AtjxR59mciYQuvs6h
MAl8S0ttMfwE1pgPmT+ixMHICsuHAM2zQ9ng/R1Vovd+6Ug5dU6pvp5U4tdJko6BE/Im/ftMmSCo
yf+5ilIlPO+8c4DmwO+lzSSBX5zCH5o2Y8lAQtYCR7ZBGVNlJS3v2KKIbsFaZvvcRVKRONK5DFIE
81y6ZlDiX/wL/MiYOJ6iH2WPCwF6RS+ShhchGytUZ4ob9JGsXwknHreyAZLpaeUuo4Qhs0tFt8Wg
E+FQ0t6n1zZPvVwbtUcvV59x2yuebhLh9jhVkt3G9mlp9soihjK8RdEdkxsJRVZ4/Id1q0/PXXvK
BtAe7PvlvdL011c8wI/57qZqqK8LyfQgX5JRogEfnoIC5JG45Qv/NAHXLDb5ghKnOr1xIb9K0dIx
+kEt9/VOEK1o2JzWsihKXDXVMu7kQaotYofHa+DoqNGbkqeBYz8LaYN+/lY+0jqfodpGdLXSqOOm
/nneJLy1lh/7jqht6P5QGU4WQj8snibZsgJ+AemEkm/bPnvMvWXHc9ylkmy9lsvP2/5zPUUnAh7g
kmQmYZd+FC913TdJFK+B9fF2WmXhrYIA8lTU8gSGxwhLo9UrPks7zhgkj+hdlnzek1ODrRGVAvCd
Ras2sB+wfivNQ93uVmgNvRDhTj3VhVpn4w2uUNaho5TG4QDcquAAA9y3NkqVuH7PRZ1GF/RkVptU
viJUJLwmch9OU8yfCj1CMlUdqtZJ4dcHTb7n5TBq3qjaVc8mN1eUuBAUgV42KxzEwPMCnaYGaK6T
c4WQ510gn/plnkt9fHFZa7r0ovzySM/NyjcgkjL/j2S1NyCbjC6+jMusCY7erQMl5sJo4eCPgKC5
w1J8fn2y+HFU88PuLp6sEgV6hf1WcEYXD+FJzqXN6227GkKPSmpPLcNJ4UEoTjNOAEu8mCQbozFf
gP+z7jjkFY7dBgp1WnA2osZMat0Y5BMVmNXy+3H3T3oqHemyPD9Q/XvQ5+G/vZLu8QFtBPkOCAJV
HwXp6deDPO806nvgHY6kBrn92iiWCmj5dSN5K5nmf5CzXuGHF6ZM1mQXVEkpGeDDPLPgZGf+JR+l
tDBDIBfT9LpGC1CI0g0mOD3IC+yY1Etai2pslbT4KCzN/B59LzKzCDVyeAdyGQzRzzKJA62wXPwi
eoU7zntZVmVaCQrafrFXXhmc6Ng7JAT7yomBHYmp0F5I0WQ6Ge6UCxmuSHzUoLzShVmCRmsYfEAT
qu1NlqafykSUXZG9PX6XoqBKnavGoOpVE6vH1DPTDhq/gs6MAJlGRe/wkwQR49lY/SQWmzJBTjRB
PMFVfNFTTLD5tmErhjtbjOJKq/S+5PiQ2hhlXrmXuNlZlL3zNLiR0Pm/Cto3DnoDlfILveapQwEh
kaNn8GDRvzS8HgcNTJGrzwNtgGrHaIC5knj6RwiTkwVARgpz5Y57EPwn6sgqRSuyvNkeduPKVbrc
EB0aQE0OxKBxTzUtRxSxtsrenonyysoLgUS8gkMzsxMZkn4nN6u+iMpA50/+9v3JCJbvcEcol2FY
/gAygruHnwl0S7L4obkIG8MESA4oKceHiepsaKAHqJOOwZQm0SEhmAdyKJDbkWJiO79m8bHCtVWm
4x9ow3NIre6LmrmDaaO6QS5kdgzA56Ylok8Sz+noRg0WniC+CwLRCVhLifAUS/L7G5QXEE8h5ZUX
9w3vqNAlQKh1azeMGMmm5s1CHf1iwjGaX02/5uU6dqJ99oSBWh7WhPqNgno0i3Jh+55dGQ49Yb5s
KUihN5hWORSbntZeueBJhpSR2ax93m/DGeQppekVCQuZk+Jxvd/r6woCsMqx9Ifl9Sx7eS1kBG67
eQAezEkhVl/D2Qi94/xa4+SH+0+jmf5klM0wOL4pgugFXCDDCTFOhTy3SLAqDKBdkx3hAWR5KP0G
zFKDjWKVcLMuj55xyNQrc5LUyMDyD4NX9jNhvQKMurco92Ic2x4K8hv8Wh5zqqL3I+gu+lnprsq1
gDGA4saA3Vw1n63lh+Fckg4NifdsYnSuAfs8Wf59k0WFNOEGVL6VmiFOUlgy1SJMiGg2vX7hWIeJ
SZ9C/ucNBonUHssS0mO0znUunsZXkhqf3mPmzxG/0Kf0pjtD5ED+gPAF3yF3SC+jHkWwB7/6ESD2
Fw5Hrbt14uHpv2St/wsvGify4yRojKWadC99rd/yHFVnNapms4fOBSQYNZbykAOE0afICF3mp0qS
oUaJczD7XvWaLWfeYNYncNNRqTMYNmDUFR9MGrG5b26EF0F4Plm7iYXInllpnkNyXVcoTM7nyme0
+Nye2fyu79IhXOIAwpAydh8I801ZBWHRIfk5tEUpio/RyEgPkJhHAY8QSgdBDq91JyaiZXFIJZG2
AH+cSq38IgToT2RwgrEHL7okgpn913J799Ot7tw6+rfScuCHReMhZyfaiHbakSmQMdPSDz867cZf
5fJ8fwf5DzCkc8czzpNlWGgx7UQYqHOa0fdsJ2SF0/UAaYjPG9cfTUFbZ98h+ppTTfastTTbh7EM
dSSI6UNW2nMLPWUABJXTg3jJhiOKJ4hhQWaSQRqtG1NnkmkhooQvjKE0rfkSRj+M4S/Odv/7/13/
ljMCO5lrLtCmFB9WNbJi2XUxvnnJ8PDYWm01g8jnCUOvldfgNeQ6vDfMIAPwGnfleX5+V5tK2sfI
t3dN/mlyxKMA/r0xj61kwHLGRywlwosEJCIwYQR446ndWoay5MScVQAbB9z39xl+XjLiHmjK4ZTS
YZOjO0iQMynwX7mu7rWgefxtZV2o4FyneLlgjIiBSBnRQ8xJhj4r5lOASs3z4hJmBD9NZfXwshcY
yC5ZbXu9w/99nrCBKbKOHWXUoLoCadv6GKu3MgUC67b/4VLbUmDgNV923f6Vs8H+0b01d6vaqHba
Ig+sOt5GTYIuiIgWAPrHKOaVougpEGF+as173ZUIXbKPMLyTdqDqSFNqFbznAigrpIRMEKyXL3CJ
EDL3/PUELbLdlincijaec4V/OlCPXnnNcj+PclE5K1jQa5tP3Wkq06q3y8vFf098ev9lGmrasdLd
16pZUCKFuhiiAst+EBDwKHnleIQdVCHeSK90JNlB01/GXfEny/kTa0VslJXQOwnHueyUF+S7IoMr
1ozYqMP2R0rXK5ly/sZAcqUNQwf8YCKgcr0DW97DmlJXCeHp7gbsGve7XkzyYWSfNITxBvnGHTdf
ypFQpARpCMg127IHRrRa/PpE+LYZlrcLVCFe5Yf39ksiOUuqS2FJ5oCNrMZm17JOreLHnp9xkvXj
e8PiopLaZzbBJbGf5uMKdJZXhVg0lKPkuNPK0soOi612Gv4p7wICkGEH6c33w3ZHltXCyzWxxpyX
Y3mURZAAk5SDdKBfi0BxtvvU3iLIY/efFjGQqZOfzBhyDBAFMPhm4pNQc6sk9m4uaI08xfu9VMIy
ClrY3UvbtHkcwUn9TXTs/WaDOonvKJ6VIJixqLcwls3ehWhF6N2nhGgxxuj0/SlbR/Ds89IGgCb5
p2nAmqcBXicPfyEdDLYYGZZH9jy49Hedoudfw1reJDaWAV3ppdo/VCJBafIuj3zQ2bpqXpWlRkv1
xpd31VC7HB4JPOJsLGqBVXFG0jjQiomDPEsDirLE2l9CtfcO/wveV4ByCMDVYteE1D5LWOGfI4e6
7s50YSn/CkO46T0GKJbffgIMpRlMAyvRWk5+8PcyWLxCdNm0YbD6me3boDvfScUBshR0fwufGfyW
jYv0zH6YRjtkZSO7+dzLZUu5jlTM1rlm2WEllz2lKGa6WZ4vCdMWuOzt+DCe3jgZezCZ2CuG4nfx
xM4hUQD5mRU1GmSOOTZSL1OsEIUpuisxaonOcvKiK/P+CdZ3VTHDythVNMMl13IEijb4ervc6QAH
kxbKQSAamsHfCjqwQ74Q6yXTYnYh15d5wxiDK4s7SXcybC99KgF86UtmJb7OIARwcZ8/Ay5l17H4
jwqbkQ3cgcHfrAjVQmEmOjkYC5Uh0rq/Cxwd4ZfKBjrgLBCG3W6ldqt7cSxnQCXtlmuuZCJ53QOX
+BXT7Em7MAp7X779gpE7gRc9vKaMO+3skWJStnk6B+v1XlRkBDMJz/5Q0upZaNziOFeBDI3Z9NtU
c2rW9oeUxnBrvepj2qaWb2Xwv0Q97rop1eBXwlReN+RP+OBLagFGlJ2n0qxJBK4AGKiNupbSYEdy
4FA2xKJOz5sUfw7rx3XB+m8DgQBrsnX1iaaU7b0eoAt2K8hEi9aN28eIrlDkW8Ix9khy0CQGfapq
VqrQm3PEJA9m+ONyYCdWrYTH8cFyDM1kVRfd/aV0tNPL4IquNMjUmG7Rd3Um6JbxkNXPquhcIvxS
CpvFAl9GrTZeh1NtopZmZUC0lDfLzbCtzLbjRh/BV5wrWCYA7J6X3DN1jxJjn+LtpYmBDvVMj/Ke
Wwpx7JJZQDrfBGLXhszO2wrcydxQW41HMLsNOW4bTvvlVXARhfxuEY+BFREdUGvBbGjmSQmoGc3r
mhtX92YKWhpFtv9+vKGLn7V5exaq96BmxmSk787D9X4CxojVTTy+OC+Ru1r9I3uXawnL5vlKqOmC
6sLp9LxF9E7fMUVuMAodFKqg0nQaMFghSLgm7AJGKFkeXLpIq8rSzU0wxBXEMAnQyJ94gGbIjuTQ
690Dn58NPRW6TXAuJpolU2CARSlquuNzOLnJkYaQztt6FkFKq3lN+7OskCZmUCstf7WH0AV/92UC
zvkfQv1GmFaWUeVd9QK+CgUw6cLCTWk18zq8tQE1U5vpSqV/APFYQoLSYPlL7KJ0Ol9og/vpMX10
0FukdUdDrReRqocptAPtmnsDCamrBQrpe5OuDn851ETuakETpdWxwaSVuwOlePz+JS6cwJ29KiCa
e2gIUFEXX3MxysAz5jISrAsJlp6Z0h+Wa8k2FeLQXiVIH/CqCYOZ5AbQwDY9tnjx1+W7REhnMS0s
xehN9DGzYyjsNgH2J06yDCvJW3zhEct04VZQbR+gKicjKrcJ1MAmLoaQ0oBX/6gKdmaCWCodMpiE
vkp93vd/8CVZZjxTzpfXUm9FvNnMnolXv2y/fhBGhdpXyc7J7hozq5w1yVZOjnHmJ/FA2LvnBG8N
UtqJ4RO5wJvNTCmllhP2M9mCAjrl1QdAKWVUuTUPSXzpmlrmHPCSVUeU9W3GR60nln46O879Qilg
cZEe15Ia6xhCGaOMXv+Xh8EgYEjdsuQqs6tp1Te/loOdZfopyzznV1cLtalK2IMTDc1CuZkYaR/I
1xHbdNxu/0oVZ4syDz9SOyC2YoB4B7ZfWcWee5GvIe+UcwcmMl/L5hbXaNvERfgZdlTzaUqQ2vU3
wwMgNnkeRi4kqyjruM16vFbYXRFH1BNi7eGrlH51GIDx5HopsZZ1vkbTRzgL+7hs4hjwUJTeOndI
YuDqEQH6nzepBJIZKnyEfYBZw53JE1PwOKEGxJpSzi5CWAuAd89iWmjK7kzWgaYeFbGs0SDmso2c
0gyBzlC2+nrZiZQBdPL4nZ2yIy16QlyAKLx8/EzXKbiPUoUCnxYpWAd8cpdlObY8UDTycML6wS7e
w5cQsPgphCFWd2Oz13Y5vPesBk/alwXGYHu63ldaZo6vrxyqWkcS8xpNPa8Ku7/n+oMC/XpvZCOX
HGtLIazXnLj+SXOeSs1WFjPbpv0VUmJgHLQqpu68neX0EhnG9Lg0++eLlkNCgc0SyybR6D2ClFL4
x9hU39IOvDhUfyEmumwaXInF4LJ4LfkPMbwf9UzILvpA9R75kp7Ft/2p+DiBfDPQ8VD/96s7+EpB
WVFCPYDbTVC1hDmtbmULtmiPf679+gFC56Pypl/kIxNdjNIvHnw5hbWJcD74wxC5zjiH+5wn0BMt
Zp1tgGxdqAIdEpYXJ0sMoCxanBaLoX5otBF8Rt5+LLDZVQ+5+MA/KZr/CesWEx4ACqhaV7b7rRG5
hwZOx7xUlAbCSeLsAdu1BvB5/iIPOLYGlI36XA7HXWwWeoHQtXuyznvmSlsqaOv91M8JLMLlNmJE
jbJxRySsYLoV+JBHUA0qshjU9P4SULd9KT+/HjxsLtYrOpfdTgZRhOjZlGTan0xLGkIBXZ3ucfUz
DeNg0qYiXQyLCqxT5seV5Jt8hxmn4E4YwBjSajWpeBfA8zEEUFXIpyiwVk44uOD9dJoOnxNPptW9
vY/9GW9KzEpQIdVsGDHJF20p0+LoXKq/Fqzrs3pKaPrgljPkpPzsy9IVHJsrlV8zMIX9j1mzKJUb
GwGB9j9HTYFHKXiHHfwriKg1tfxyQ9028SWTWicbH8ONJzgr/lhxIXlUtD2mC/wYurzwH1pxC6Ch
V1GcAjieJNf3+QUkWVWlAhJOUF7ZhlIRIkb7H2EKsxZLq/YFxZhFNRDoDry8mAYfFgRjX3QAsHsB
pGlkqrFlK7a+1vXr08PiQpplK9q6J6kpDnJFDl4rqe8yroTlpGWO7zRMRhDapFUAeEWYW+4kmYBJ
HyW+NUmWEopZakxBiEmH9sVh/q9D3kHTfRMQzRPm82UBApqRuAatX8noJtd+JoRE+x00a6bFUZ4V
fwI2AUfTcHTOQCL6YvfiuHLiyMTrSW9mR5Mq2lmAuf0jrm9o3GPaVDAitbIU0WMXpsR6nqJzqYCK
0JcPSEXcsDTRD0J5/Zh9QNBN5KHyDdUj+KUOxBo7YrskAcRINga5F344Ho892a7dLFiCB4aC1NKP
W2g3BiFlSl0MFJ6F6RcH5Fh7m1830yjlXNrY2Bqbkdxaqbx4Vu5swgM2dGc17ZW7YezKAMEodWv9
a21JT7xR1gmNfN7MCe1HJxu0cai+1bNbpnhWBDh2C2I1BkF6PECtX+yYKQ5K5DLLt0f524R4A8tJ
cLYWmB+B259kkVTOyiovccwVeZqmqQCABvFuxsxMEj2pUQcAqEsCTOvQVpdhS7sBbGQHyKg4HLT9
APv77c/RckUvAV+sP7jrjc2Cdik5O/vS8sR1c79OgiiqifyV976pilckofU9UaTW2+SMa6oAnheQ
wVOAONmbrxy7rj1nWYAEQigL7r6GCCmggCIcpxRB0+uVvYhOuphCQ6EnX330jxVOoL7tgHAi+Akn
HZjQ0mmngAH41ViPpy3Vt2Grt/6eZ27mWtY/JYIjPYYKRUuXDbgx24aBV5UK5Q3ttY5W6RsPdOKB
k8Gw/HiTfhdUDvZhFbSydZdRNlSeVDG4LFqNcJ6Q7TdURkS7fud2ekA4ly/rsw/HA3TIOMB0gqJw
dCUmHPhk7Ah12ytyZVwpBxLCJL4RgblIr0pWBhxk9CnBuPH7CxzKqrRepbreG3pAwNosdCadCGeJ
Wu1nD0uMzJ3LmWoL7JzwnToLZqU0O/72exr/zZSocBXjPnghd83f0bbL7peoBRx8RUSigarxmhv7
oHqnOXtoqLRp9aU+QFcUzlc1zeZxU7XDylUMB8WlhKE30qZZxNyaD9Zx494HCWup4qVhpcxvyyuX
qXRKAa6iXXTLhWMEY8Wne9XZJWMhZvypTCaFlgyl7nxAQCH8EasOgGbb6owu4JVQ70pZpHIhKmBR
rF2+TfyWONt+XJGUvOIMVY695drmcJ+igybR0A56TPb91kjGxBjuF84QDsgPXXQuOdWnrLARWIgr
JY7XxC7gdzJI7ydTSirRMl1N4qIBxLBEgUIqifRKfnPkQXXdy1cIYf1KV8xzR6cPsJr73sGcXcl9
onsrp3QVbjm/732jbKj919NdeWGO9XtXTAfSclYD5Dmut20e9qQUTeXJka1ZLKpg+N/jLLB92Y0t
ZtFByAcWF4kq3HbQburCWsx+IWny50KD9nbop5kKe3uWS/n9RmdDA49JHh7wIJufVVd1QZ2fDPj+
Wspm92H9dg6LQ8CxFZy1QOhrST80xLAXd7NO0cbMKwQGNgYp98Ms8XFBIgqW9EGR7rzDerBRynFt
ISdeM2CosVg1eu6DTNP3U6ZoX7BZe+Z/mt2VGBKQrueC2z6KdzfYmgnHF1FaUsI2Io3RRpzkw+EK
ZJ0OSWUeLdjq5oESY3h/P8yL+rmojhMM2+3V24B/ROZuBGj3DF32phHDwofbzJxCZETuRXFA0SKu
Y40KkAff+Ml/6e1xJx82f/Z+6KTgLmtqd8ZLMJxJnYPE3NuPleF9l37IUMVyfc8kDcFO+ywI0oQJ
3WKhwtOlPrmGx8V4SL4PO/xi/IX8O+7NVzPChWMp5wWU7MKgqf/BN+689DYkqbEebhe/vulPxxF1
eODDLemUANlbFaEKbQ7TKAYxBbgBC29k7yMInFGRPefkLQ+Gw6lgjLXikGdDDxKHUYtrf75tR12v
gVblaocP7p0ry//9cR1zoMrN8VXxl22xgSHw9P+qzh0DyVGcbW0yxX+57JIYalw+0YUxxIsYu5FK
2IOSfsniav22eeGYpwY9RLS+LlGO0bWvuV71tszYX/WjfZV5tKBNi5HkBDOYKUxMMseXrt+GazHi
Qj2axKCpCcysAGPpYqO5qAJCQbzHeFoFdDB22NZM7kBVitBBZBWky0Mmt1jgz2dVKmwP/v7Z6hrf
BhwSJL0YvTvT7xZcJlwRpU31aEl4Sr2hH1ugEbGjEuHKAufQ+HIXHN1ESKXNHncWsTfozJ+BYPkA
HaTRHtEmbWxCEVFMxxJMZYujR4Lvvs7nDYmFGUnaYL86v62ZrOOAsoMhg/leqA7Z2NKXUSzt3+RS
YnxTJ6tZffiSX3n7DVw4JPYwauTNn7V9kNPougdTH9GF6JWaODxqGHhAIwTZVnm4fAe4vUiUDcm1
30Y+76P4hMHHLKDmE8aRUWLe5Q5W1ImpC8q7Sz0ULyLTd3IgUYxxZJr2QTMCHqldF1+V9zkrJynn
Tarb4koHNaipJWq4b3bBMfRxULUQGsZIbu2q0BcJ0GZl/x0KhIRB7Z1vCWW4vWdRyO4P9YoX2SNA
s603kmFzj2I7TAcx5XFWQEgK4BVds8MRJix1Qm+QO3xzHc+vTKxh2oRX+rU8EnJieRXz5K6hEwu4
LQ4XzwRtKLTeV9f/nbgI5S/VevoOWgyFcgzCdeYA3FQzsgnb/aaVkwfCH55gcr6lazjBHQmae3oB
j0HeEBRWJmhG99pDYc3n7dQouzO8VNLz25aEZePrRtvLfYtCr7cO88ggWVM6gUmXZGh8cGzLax1u
/9RfKuKbkJ3USdIXa+Kq+RVTHFWr9jpPq7ZCFE+Do2HsXRvHredua6RSVsOaOGQoQwKUdKWxfhVT
KvxOD6InR8tPlWiJhZOnnbaIMeaXNBquq67uc+zTbWHN2gYcuQfXnxOs0+Bvpp6rBANO4n8XPEin
lvmTEkONX0deDx9g+ksB8eKM3DpgCQmtcZ1ZrHbOp3BS5p4wCjz4RAZIiI7PM0XgkoA1Z6S7p7vZ
DPTwm89wSam2vAAg3AyBxv7wXORvmrdX9WeCcym5S1aE6MMnl/ex+BUMSrc59GcG/oZ7BEDvMaiv
tXxWjb3EutBowRetBUX5BivZxyYTiF+4EzIp43NaSmKffSsNTiwGW41E03XZKM1B6ZNgIQ9BGtVJ
TaQVAd7iJp73cGWXeO/o/dMW1RBVFlan6IEljMpgHECLqSlvQPqHOctnS2IGop6+je77jB5aCCMO
Do+ooWvsKxML3Xs9zqWNAZX5znax/w5pVowSUcfnFCChVwpuwpNN+w6/aDbs8hM6RsGCOzwUdvmi
pCOJNBrOm5bqHYujD3TWrQmsjB+tIr5RMKuayEE3CxNEfqmV4X/nHXXiDe2IlX6i5Lwhz2re74wt
aUF7Aw2jsOVOUYDCOrvPbSKvlu8PunxQpJhM2JqN5SaAt2rzZIklZRfjvM9nbxk2E5ZMuIlrDdB3
9K70BtjnXUZcdq5SbBXnGn35U1+MQvFdD2z3gaz6iAg8q8DKpFrxn6BelkaUJSWUYQfv1ebcQxZe
QzpJ/v/4pDkWS0nmuQRmr8ZhtGYlj7olzAqCNd9L8fNPUbeDsrFqsGWUjZq0DhzIY+QJcBgb7V8a
JFPBI42spZLj6D1bnIx/nORmi57trEKVmunkuclrtiKx/1zKNiGv+y5+/QBPaj0hSiMlUGOtIIaX
jnk5Aa43ZuEVSPl+0Htv4i50rxk8YtiRRr8QuRHJ8QghlmjXME29UIzNT+HtoOoXJiks+WWXNbJg
NHGPfjQdWGdeQiuTWkAIxsCXWLt4cvAuqPlbTp4ayNi2hzQ0ZI2p2w4WwcWYJxCL3aHK4YuXrGec
Jtabqv6/Xp9sfrc/8Zo528dyY5Nohyx40jdghmxrXSSgOSccZ2POg9PaIPe0tZZCfaXZ4g5nGhzm
DT+1ueqQ5H2ZpMQpS04E3D+A7FqANqx0DQsJ40IVYLPitfZlzvvTVcv6hhKWIV4maT3OZdPpcZkZ
Bizp69m8dYD21cvH2g/chcEAYoU8T1Z5ezmh0aoGIxHc4aKbSvFe8OC7OBvrLxMabfhIXedHQR8v
YGmvq5T1bBC6U17HHIApJ/AoJyHp5I+spMITbBeFcRfzcsbL9ilAKrFtItL/alpdafIP0Tb55r0g
JvWhGLXaDWO0unXkFuuAzeZw07gCcfHClG3xQMNwVnV8WX2iSa5xoywPzuHWjanFoiNe9V5PMcUK
0Aa4w3Spzdit4aUIyZHf8mAC5XuVSQMHors5MU7Wxdlu8UFsOIWEffRNQ1MOq2nbIaxvrryaFDfU
F+JovT6OHwjJqU9Ml97uucm4T4mYWr42PN5WbTSDqY8rsT4xv49XRIpIccefxaR1inoKwizUO8OZ
jzE6iG74cUplYK3I1Q92Yu4osmkVqYfTQENve5Ps45uKOeEdzbo/h9H82b9KGDn9lSVzO2kcZIPE
HSZdcVKVpmgI7unfPYvyefo2RQJivc+HMEkcPho/9ryS3sP1Oz4oHRRIMa65xKvHrkm+zgAUcwtB
qx6tUYJnZnA6Qje0OkWWT+1rzcMrBoHU/GT0LTKdgBsyDW9CdQXw4tHcGJ+tpX1TzbQ68W7crZaS
vR0jz/SHf5VlYjZWRLArw1d+KeweganlhP0WIiOyK9jDCINT59YFzTE14n6twB3eUpp5maxXHFvL
tBPjoL05MaX/27zafPWQOGikjhuy9s4/r/pcszziLI6bjXMlkFZ3Ldy6h1nmhnYKbj7uDU+EDePX
eQ==
`pragma protect end_protected
