`define module_name I2C_MASTER_Top
