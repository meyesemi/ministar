// ===========Oooo==========================================Oooo========
// =  Copyright (C) 2014-2020 Shandong Gowin Semiconductor Technology Co.,Ltd.
// =                     All rights reserved.
// =====================================================================
//
//  __      __      __
//  \ \    /  \    / /   [File name   ] ROM549x17.v
//   \ \  / /\ \  / /    [Description ] Verilog file for the DPHY testbench design
//    \ \/ /  \ \/ /     [Timestamp   ] Tue Mar 24 15:30:00 2020
//     \  /    \  /      [version     ] 1.0
//      \/      \/
// --------------------------------------------------------------------
// Code Revision History :
// --------------------------------------------------------------------
// Ver: | Author |Mod. Date |Changes Made:
// V1.0 | XX     |24/03/20  |Initial version
// ===========Oooo==========================================Oooo========
`timescale 1ns/1ps

module ROM549x17(
    clk   ,
    rstn  ,
    dout  
    );

  input         clk   ;
  input         rstn  ;
  output [16:0] dout  ;

  reg    [16:0] dout  ;
  reg     [9:0] addr  ;

  always@(posedge clk or negedge rstn)
  begin
    if(!rstn)
      addr <= 'b0;
    else
      addr <= addr + 1'b1;
  end

  always@(posedge clk)
  begin
    case(addr)
      0   :   dout <= 17'h00000;     
      1	  :   dout <= 17'h00000;     
      2	  :   dout <= 17'h00000;     
      3	  :   dout <= 17'h00000;     
      4	  :   dout <= 17'h00000;     
      5	  :   dout <= 17'h00000;     
      6	  :   dout <= 17'h00000;     
      7	  :   dout <= 17'h00000;     
      8	  :   dout <= 17'h00000;     
      9	  :   dout <= 17'h00000;     
      10	:   dout <= 17'h00000;     
      11	:   dout <= 17'h00000;     
      12	:   dout <= 17'h00000;     
      13	:   dout <= 17'h00000;     
      14	:   dout <= 17'h00000;     
      15	:   dout <= 17'h00000;     
      16	:   dout <= 17'h00000;     
      17	:   dout <= 17'h00000;     
      18	:   dout <= 17'h00000;     
      19	:   dout <= 17'h00000;     
      20	:   dout <= 17'h00000;     
      21	:   dout <= 17'h00000;     
      22	:   dout <= 17'h00000;     
      23	:   dout <= 17'h00000;     
      24	:   dout <= 17'h00000;     
      25	:   dout <= 17'h00000;     
      26	:   dout <= 17'h00000;     
      27	:   dout <= 17'h00000;     
      28	:   dout <= 17'h00000;     
      29	:   dout <= 17'h00000;     
      30	:   dout <= 17'h00000;     
      31	:   dout <= 17'h00000;     
      32	:   dout <= 17'h00000;     
      33	:   dout <= 17'h00000;     
      34	:   dout <= 17'h00000;     
      35	:   dout <= 17'h00000;     
      36	:   dout <= 17'h00000;     
      37	:   dout <= 17'h00000;     
      38	:   dout <= 17'h00000;     
      39	:   dout <= 17'h00000;     
      40	:   dout <= 17'h00000;     
      41	:   dout <= 17'h00000;     
      42	:   dout <= 17'h00000;     
      43	:   dout <= 17'h00000;     
      44	:   dout <= 17'h00000;     
      45	:   dout <= 17'h00000;     
      46	:   dout <= 17'h00000;     
      47	:   dout <= 17'h00000;     
      48	:   dout <= 17'h00000;     
      49	:   dout <= 17'h00000;     
      50	:   dout <= 17'h00000;     
      51	:   dout <= 17'h00000;     
      52	:   dout <= 17'h00000;     
      53	:   dout <= 17'h00000;     
      54	:   dout <= 17'h00000;     
      55	:   dout <= 17'h00000;     
      56	:   dout <= 17'h00000;     
      57	:   dout <= 17'h00000;     
      58	:   dout <= 17'h00000;     
      59	:   dout <= 17'h10000;     
      60	:   dout <= 17'h10000;     
      61	:   dout <= 17'h10000;     
      62	:   dout <= 17'h10000;     
      63	:   dout <= 17'h10000;     
      64	:   dout <= 17'h10000;     
      65	:   dout <= 17'h137b8;     
      66	:   dout <= 17'h12a2a;     
      67	:   dout <= 17'h10000;     
      68	:   dout <= 17'h18080;     
      69	:   dout <= 17'h14040;     
      70	:   dout <= 17'h1c0c0;     
      71	:   dout <= 17'h12020;     
      72	:   dout <= 17'h1a0a0;     
      73	:   dout <= 17'h16060;     
      74	:   dout <= 17'h1e0e0;     
      75	:   dout <= 17'h10000;     
      76	:   dout <= 17'h18080;     
      77	:   dout <= 17'h14040;     
      78	:   dout <= 17'h1c0c0;     
      79	:   dout <= 17'h12020;     
      80	:   dout <= 17'h1a0a0;     
      81	:   dout <= 17'h16060;     
      82	:   dout <= 17'h1e0e0;     
      83	:   dout <= 17'h10000;     
      84	:   dout <= 17'h18080;     
      85	:   dout <= 17'h14040;     
      86	:   dout <= 17'h1c0c0;     
      87	:   dout <= 17'h12020;     
      88	:   dout <= 17'h1a0a0;     
      89	:   dout <= 17'h16060;     
      90	:   dout <= 17'h1e0e0;     
      91	:   dout <= 17'h10000;     
      92	:   dout <= 17'h18080;     
      93	:   dout <= 17'h14040;     
      94	:   dout <= 17'h1c0c0;     
      95	:   dout <= 17'h12020;     
      96	:   dout <= 17'h1a0a0;     
      97	:   dout <= 17'h16060;     
      98	:   dout <= 17'h1e0e0;     
      99	:   dout <= 17'h10000;     
      100	:   dout <= 17'h18080;     
      101	:   dout <= 17'h14040;     
      102	:   dout <= 17'h1c0c0;     
      103	:   dout <= 17'h12020;     
      104	:   dout <= 17'h1a0a0;     
      105	:   dout <= 17'h16060;     
      106	:   dout <= 17'h1e0e0;     
      107	:   dout <= 17'h10000;     
      108	:   dout <= 17'h18080;     
      109	:   dout <= 17'h14040;     
      110	:   dout <= 17'h1c0c0;     
      111	:   dout <= 17'h12020;     
      112	:   dout <= 17'h1a0a0;     
      113	:   dout <= 17'h16060;     
      114	:   dout <= 17'h1e0e0;     
      115	:   dout <= 17'h10000;     
      116	:   dout <= 17'h18080;     
      117	:   dout <= 17'h14040;     
      118	:   dout <= 17'h1c0c0;     
      119	:   dout <= 17'h12020;     
      120	:   dout <= 17'h1a0a0;     
      121	:   dout <= 17'h16060;     
      122	:   dout <= 17'h1e0e0;     
      123	:   dout <= 17'h10000;     
      124	:   dout <= 17'h18080;     
      125	:   dout <= 17'h14040;     
      126	:   dout <= 17'h1c0c0;     
      127	:   dout <= 17'h12020;     
      128	:   dout <= 17'h1a0a0;     
      129	:   dout <= 17'h16060;     
      130	:   dout <= 17'h1e0e0;     
      131	:   dout <= 17'h10000;     
      132	:   dout <= 17'h18080;     
      133	:   dout <= 17'h14040;     
      134	:   dout <= 17'h1c0c0;     
      135	:   dout <= 17'h12020;     
      136	:   dout <= 17'h1a0a0;     
      137	:   dout <= 17'h16060;     
      138	:   dout <= 17'h1e0e0;     
      139	:   dout <= 17'h10000;     
      140	:   dout <= 17'h18080;     
      141	:   dout <= 17'h14040;     
      142	:   dout <= 17'h1c0c0;     
      143	:   dout <= 17'h12020;     
      144	:   dout <= 17'h1a0a0;     
      145	:   dout <= 17'h16060;     
      146	:   dout <= 17'h1e0e0;     
      147	:   dout <= 17'h10000;     
      148	:   dout <= 17'h18080;     
      149	:   dout <= 17'h14040;     
      150	:   dout <= 17'h1c0c0;     
      151	:   dout <= 17'h12020;     
      152	:   dout <= 17'h1a0a0;     
      153	:   dout <= 17'h16060;     
      154	:   dout <= 17'h1e0e0;     
      155	:   dout <= 17'h10000;     
      156	:   dout <= 17'h18080;     
      157	:   dout <= 17'h14040;     
      158	:   dout <= 17'h1c0c0;     
      159	:   dout <= 17'h12020;     
      160	:   dout <= 17'h1a0a0;     
      161	:   dout <= 17'h16060;     
      162	:   dout <= 17'h1e0e0;     
      163	:   dout <= 17'h10000;     
      164	:   dout <= 17'h18080;     
      165	:   dout <= 17'h14040;     
      166	:   dout <= 17'h1c0c0;     
      167	:   dout <= 17'h12020;     
      168	:   dout <= 17'h1a0a0;     
      169	:   dout <= 17'h16060;     
      170	:   dout <= 17'h1e0e0;     
      171	:   dout <= 17'h10000;     
      172	:   dout <= 17'h18080;     
      173	:   dout <= 17'h14040;     
      174	:   dout <= 17'h1c0c0;     
      175	:   dout <= 17'h12020;     
      176	:   dout <= 17'h1a0a0;     
      177	:   dout <= 17'h16060;     
      178	:   dout <= 17'h1e0e0;     
      179	:   dout <= 17'h10000;     
      180	:   dout <= 17'h18080;     
      181	:   dout <= 17'h14040;     
      182	:   dout <= 17'h1c0c0;     
      183	:   dout <= 17'h12020;     
      184	:   dout <= 17'h1a0a0;     
      185	:   dout <= 17'h16060;     
      186	:   dout <= 17'h1e0e0;     
      187	:   dout <= 17'h10000;     
      188	:   dout <= 17'h18080;     
      189	:   dout <= 17'h14040;     
      190	:   dout <= 17'h1c0c0;     
      191	:   dout <= 17'h12020;     
      192	:   dout <= 17'h1a0a0;     
      193	:   dout <= 17'h16060;     
      194	:   dout <= 17'h1e0e0;     
      195	:   dout <= 17'h10000;     
      196	:   dout <= 17'h18080;     
      197	:   dout <= 17'h14040;     
      198	:   dout <= 17'h1c0c0;     
      199	:   dout <= 17'h12020;     
      200	:   dout <= 17'h1a0a0;     
      201	:   dout <= 17'h16060;     
      202	:   dout <= 17'h1e0e0;     
      203	:   dout <= 17'h10000;     
      204	:   dout <= 17'h18080;     
      205	:   dout <= 17'h14040;     
      206	:   dout <= 17'h1c0c0;     
      207	:   dout <= 17'h12020;     
      208	:   dout <= 17'h1a0a0;     
      209	:   dout <= 17'h16060;     
      210	:   dout <= 17'h1e0e0;     
      211	:   dout <= 17'h10000;     
      212	:   dout <= 17'h18080;     
      213	:   dout <= 17'h14040;     
      214	:   dout <= 17'h1c0c0;     
      215	:   dout <= 17'h12020;     
      216	:   dout <= 17'h1a0a0;     
      217	:   dout <= 17'h16060;     
      218	:   dout <= 17'h1e0e0;     
      219	:   dout <= 17'h10000;     
      220	:   dout <= 17'h18080;     
      221	:   dout <= 17'h14040;     
      222	:   dout <= 17'h1c0c0;     
      223	:   dout <= 17'h12020;     
      224	:   dout <= 17'h1a0a0;     
      225	:   dout <= 17'h16060;     
      226	:   dout <= 17'h1e0e0;     
      227	:   dout <= 17'h10000;     
      228	:   dout <= 17'h18080;     
      229	:   dout <= 17'h14040;     
      230	:   dout <= 17'h1c0c0;     
      231	:   dout <= 17'h12020;     
      232	:   dout <= 17'h1a0a0;     
      233	:   dout <= 17'h16060;     
      234	:   dout <= 17'h1e0e0;     
      235	:   dout <= 17'h10000;     
      236	:   dout <= 17'h18080;     
      237	:   dout <= 17'h14040;     
      238	:   dout <= 17'h1c0c0;     
      239	:   dout <= 17'h12020;     
      240	:   dout <= 17'h1a0a0;     
      241	:   dout <= 17'h16060;     
      242	:   dout <= 17'h1e0e0;     
      243	:   dout <= 17'h10000;     
      244	:   dout <= 17'h18080;     
      245	:   dout <= 17'h14040;     
      246	:   dout <= 17'h1c0c0;     
      247	:   dout <= 17'h12020;     
      248	:   dout <= 17'h1a0a0;     
      249	:   dout <= 17'h16060;     
      250	:   dout <= 17'h1e0e0;     
      251	:   dout <= 17'h10000;     
      252	:   dout <= 17'h18080;     
      253	:   dout <= 17'h14040;     
      254	:   dout <= 17'h1c0c0;     
      255	:   dout <= 17'h12020;     
      256	:   dout <= 17'h1a0a0;     
      257	:   dout <= 17'h16060;     
      258	:   dout <= 17'h1e0e0;     
      259	:   dout <= 17'h10000;     
      260	:   dout <= 17'h18080;     
      261	:   dout <= 17'h14040;     
      262	:   dout <= 17'h1c0c0;     
      263	:   dout <= 17'h12020;     
      264	:   dout <= 17'h1a0a0;     
      265	:   dout <= 17'h16060;     
      266	:   dout <= 17'h1e0e0;     
      267	:   dout <= 17'h10000;     
      268	:   dout <= 17'h18080;     
      269	:   dout <= 17'h14040;     
      270	:   dout <= 17'h1c0c0;     
      271	:   dout <= 17'h12020;     
      272	:   dout <= 17'h1a0a0;     
      273	:   dout <= 17'h16060;     
      274	:   dout <= 17'h1e0e0;     
      275	:   dout <= 17'h10000;     
      276	:   dout <= 17'h18080;     
      277	:   dout <= 17'h14040;     
      278	:   dout <= 17'h1c0c0;     
      279	:   dout <= 17'h12020;     
      280	:   dout <= 17'h1a0a0;     
      281	:   dout <= 17'h16060;     
      282	:   dout <= 17'h1e0e0;     
      283	:   dout <= 17'h10000;     
      284	:   dout <= 17'h18080;     
      285	:   dout <= 17'h14040;     
      286	:   dout <= 17'h1c0c0;     
      287	:   dout <= 17'h12020;     
      288	:   dout <= 17'h1a0a0;     
      289	:   dout <= 17'h16060;     
      290	:   dout <= 17'h1e0e0;     
      291	:   dout <= 17'h10000;     
      292	:   dout <= 17'h18080;     
      293	:   dout <= 17'h14040;     
      294	:   dout <= 17'h1c0c0;     
      295	:   dout <= 17'h12020;     
      296	:   dout <= 17'h1a0a0;     
      297	:   dout <= 17'h16060;     
      298	:   dout <= 17'h1e0e0;     
      299	:   dout <= 17'h10000;     
      300	:   dout <= 17'h18080;     
      301	:   dout <= 17'h14040;     
      302	:   dout <= 17'h1c0c0;     
      303	:   dout <= 17'h12020;     
      304	:   dout <= 17'h1a0a0;     
      305	:   dout <= 17'h16060;     
      306	:   dout <= 17'h1e0e0;     
      307	:   dout <= 17'h10000;     
      308	:   dout <= 17'h18080;     
      309	:   dout <= 17'h14040;     
      310	:   dout <= 17'h1c0c0;     
      311	:   dout <= 17'h12020;     
      312	:   dout <= 17'h1a0a0;     
      313	:   dout <= 17'h16060;     
      314	:   dout <= 17'h1e0e0;     
      315	:   dout <= 17'h10000;     
      316	:   dout <= 17'h18080;     
      317	:   dout <= 17'h14040;     
      318	:   dout <= 17'h1c0c0;     
      319	:   dout <= 17'h12020;     
      320	:   dout <= 17'h1a0a0;     
      321	:   dout <= 17'h16060;     
      322	:   dout <= 17'h1e0e0;     
      323	:   dout <= 17'h10000;     
      324	:   dout <= 17'h18080;     
      325	:   dout <= 17'h14040;     
      326	:   dout <= 17'h1c0c0;     
      327	:   dout <= 17'h12020;     
      328	:   dout <= 17'h1a0a0;     
      329	:   dout <= 17'h16060;     
      330	:   dout <= 17'h1e0e0;     
      331	:   dout <= 17'h10000;     
      332	:   dout <= 17'h18080;     
      333	:   dout <= 17'h14040;     
      334	:   dout <= 17'h1c0c0;     
      335	:   dout <= 17'h12020;     
      336	:   dout <= 17'h1a0a0;     
      337	:   dout <= 17'h16060;     
      338	:   dout <= 17'h1e0e0;     
      339	:   dout <= 17'h10000;     
      340	:   dout <= 17'h18080;     
      341	:   dout <= 17'h14040;     
      342	:   dout <= 17'h1c0c0;     
      343	:   dout <= 17'h12020;     
      344	:   dout <= 17'h1a0a0;     
      345	:   dout <= 17'h16060;     
      346	:   dout <= 17'h1e0e0;     
      347	:   dout <= 17'h10000;     
      348	:   dout <= 17'h18080;     
      349	:   dout <= 17'h14040;     
      350	:   dout <= 17'h1c0c0;     
      351	:   dout <= 17'h12020;     
      352	:   dout <= 17'h1a0a0;     
      353	:   dout <= 17'h16060;     
      354	:   dout <= 17'h1e0e0;     
      355	:   dout <= 17'h10000;     
      356	:   dout <= 17'h18080;     
      357	:   dout <= 17'h14040;     
      358	:   dout <= 17'h1c0c0;     
      359	:   dout <= 17'h12020;     
      360	:   dout <= 17'h1a0a0;     
      361	:   dout <= 17'h16060;     
      362	:   dout <= 17'h1e0e0;     
      363	:   dout <= 17'h10000;     
      364	:   dout <= 17'h18080;     
      365	:   dout <= 17'h14040;     
      366	:   dout <= 17'h1c0c0;     
      367	:   dout <= 17'h12020;     
      368	:   dout <= 17'h1a0a0;     
      369	:   dout <= 17'h16060;     
      370	:   dout <= 17'h1e0e0;     
      371	:   dout <= 17'h10000;     
      372	:   dout <= 17'h18080;     
      373	:   dout <= 17'h14040;     
      374	:   dout <= 17'h1c0c0;     
      375	:   dout <= 17'h12020;     
      376	:   dout <= 17'h1a0a0;     
      377	:   dout <= 17'h16060;     
      378	:   dout <= 17'h1e0e0;     
      379	:   dout <= 17'h10000;     
      380	:   dout <= 17'h18080;     
      381	:   dout <= 17'h14040;     
      382	:   dout <= 17'h1c0c0;     
      383	:   dout <= 17'h12020;     
      384	:   dout <= 17'h1a0a0;     
      385	:   dout <= 17'h16060;     
      386	:   dout <= 17'h1e0e0;     
      387	:   dout <= 17'h10000;     
      388	:   dout <= 17'h18080;     
      389	:   dout <= 17'h14040;     
      390	:   dout <= 17'h1c0c0;     
      391	:   dout <= 17'h12020;     
      392	:   dout <= 17'h1a0a0;     
      393	:   dout <= 17'h16060;     
      394	:   dout <= 17'h1e0e0;     
      395	:   dout <= 17'h10000;     
      396	:   dout <= 17'h18080;     
      397	:   dout <= 17'h14040;     
      398	:   dout <= 17'h1c0c0;     
      399	:   dout <= 17'h12020;     
      400	:   dout <= 17'h1a0a0;     
      401	:   dout <= 17'h16060;     
      402	:   dout <= 17'h1e0e0;     
      403	:   dout <= 17'h10000;     
      404	:   dout <= 17'h18080;     
      405	:   dout <= 17'h14040;     
      406	:   dout <= 17'h1c0c0;     
      407	:   dout <= 17'h12020;     
      408	:   dout <= 17'h1a0a0;     
      409	:   dout <= 17'h16060;     
      410	:   dout <= 17'h1e0e0;     
      411	:   dout <= 17'h10000;     
      412	:   dout <= 17'h18080;     
      413	:   dout <= 17'h14040;     
      414	:   dout <= 17'h1c0c0;     
      415	:   dout <= 17'h12020;     
      416	:   dout <= 17'h1a0a0;     
      417	:   dout <= 17'h16060;     
      418	:   dout <= 17'h1e0e0;     
      419	:   dout <= 17'h10000;     
      420	:   dout <= 17'h18080;     
      421	:   dout <= 17'h14040;     
      422	:   dout <= 17'h1c0c0;     
      423	:   dout <= 17'h12020;     
      424	:   dout <= 17'h1a0a0;     
      425	:   dout <= 17'h16060;     
      426	:   dout <= 17'h1e0e0;     
      427	:   dout <= 17'h10000;     
      428	:   dout <= 17'h18080;     
      429	:   dout <= 17'h14040;     
      430	:   dout <= 17'h1c0c0;     
      431	:   dout <= 17'h12020;     
      432	:   dout <= 17'h1a0a0;     
      433	:   dout <= 17'h16060;     
      434	:   dout <= 17'h1e0e0;     
      435	:   dout <= 17'h10000;     
      436	:   dout <= 17'h18080;     
      437	:   dout <= 17'h14040;     
      438	:   dout <= 17'h1c0c0;     
      439	:   dout <= 17'h12020;     
      440	:   dout <= 17'h1a0a0;     
      441	:   dout <= 17'h16060;     
      442	:   dout <= 17'h1e0e0;     
      443	:   dout <= 17'h10000;     
      444	:   dout <= 17'h18080;     
      445	:   dout <= 17'h14040;     
      446	:   dout <= 17'h1c0c0;     
      447	:   dout <= 17'h12020;     
      448	:   dout <= 17'h1a0a0;     
      449	:   dout <= 17'h16060;     
      450	:   dout <= 17'h1e0e0;     
      451	:   dout <= 17'h10000;     
      452	:   dout <= 17'h18080;     
      453	:   dout <= 17'h14040;     
      454	:   dout <= 17'h1c0c0;     
      455	:   dout <= 17'h12020;     
      456	:   dout <= 17'h1a0a0;     
      457	:   dout <= 17'h16060;     
      458	:   dout <= 17'h1e0e0;     
      459	:   dout <= 17'h10000;     
      460	:   dout <= 17'h18080;     
      461	:   dout <= 17'h14040;     
      462	:   dout <= 17'h1c0c0;     
      463	:   dout <= 17'h12020;     
      464	:   dout <= 17'h1a0a0;     
      465	:   dout <= 17'h16060;     
      466	:   dout <= 17'h1e0e0;     
      467	:   dout <= 17'h10000;     
      468	:   dout <= 17'h18080;     
      469	:   dout <= 17'h14040;     
      470	:   dout <= 17'h1c0c0;     
      471	:   dout <= 17'h12020;     
      472	:   dout <= 17'h1a0a0;     
      473	:   dout <= 17'h16060;     
      474	:   dout <= 17'h1e0e0;     
      475	:   dout <= 17'h10000;     
      476	:   dout <= 17'h18080;     
      477	:   dout <= 17'h14040;     
      478	:   dout <= 17'h1c0c0;     
      479	:   dout <= 17'h12020;     
      480	:   dout <= 17'h1a0a0;     
      481	:   dout <= 17'h16060;     
      482	:   dout <= 17'h1e0e0;     
      483	:   dout <= 17'h10000;     
      484	:   dout <= 17'h18080;     
      485	:   dout <= 17'h14040;     
      486	:   dout <= 17'h1c0c0;     
      487	:   dout <= 17'h12020;     
      488	:   dout <= 17'h1a0a0;     
      489	:   dout <= 17'h16060;     
      490	:   dout <= 17'h1e0e0;     
      491	:   dout <= 17'h10000;     
      492	:   dout <= 17'h18080;     
      493	:   dout <= 17'h14040;     
      494	:   dout <= 17'h1c0c0;     
      495	:   dout <= 17'h12020;     
      496	:   dout <= 17'h1a0a0;     
      497	:   dout <= 17'h16060;     
      498	:   dout <= 17'h1e0e0;     
      499	:   dout <= 17'h10000;     
      500	:   dout <= 17'h18080;     
      501	:   dout <= 17'h14040;     
      502	:   dout <= 17'h1c0c0;     
      503	:   dout <= 17'h12020;     
      504	:   dout <= 17'h1a0a0;     
      505	:   dout <= 17'h16060;     
      506	:   dout <= 17'h1e0e0;     
      507	:   dout <= 17'h10000;     
      508	:   dout <= 17'h18080;     
      509	:   dout <= 17'h14040;     
      510	:   dout <= 17'h1c0c0;     
      511	:   dout <= 17'h12020;     
      512	:   dout <= 17'h1a0a0;     
      513	:   dout <= 17'h16060;     
      514	:   dout <= 17'h1e0e0;     
      515	:   dout <= 17'h10000;     
      516	:   dout <= 17'h18080;     
      517	:   dout <= 17'h14040;     
      518	:   dout <= 17'h1c0c0;     
      519	:   dout <= 17'h12020;     
      520	:   dout <= 17'h1a0a0;     
      521	:   dout <= 17'h16060;     
      522	:   dout <= 17'h1e0e0;     
      523	:   dout <= 17'h10000;     
      524	:   dout <= 17'h18080;     
      525	:   dout <= 17'h14040;     
      526	:   dout <= 17'h1c0c0;     
      527	:   dout <= 17'h12020;     
      528	:   dout <= 17'h1a0a0;     
      529	:   dout <= 17'h16060;     
      530	:   dout <= 17'h1e0e0;     
      531	:   dout <= 17'h10000;     
      532	:   dout <= 17'h18080;     
      533	:   dout <= 17'h14040;     
      534	:   dout <= 17'h1c0c0;     
      535	:   dout <= 17'h12020;     
      536	:   dout <= 17'h1a0a0;     
      537	:   dout <= 17'h16060;     
      538	:   dout <= 17'h1e0e0;     
      539	:   dout <= 17'h10000;     
      540	:   dout <= 17'h18080;     
      541	:   dout <= 17'h14040;     
      542	:   dout <= 17'h1c0c0;     
      543	:   dout <= 17'h12020;     
      544	:   dout <= 17'h1a0a0;     
      545	:   dout <= 17'h16060;     
      546	:   dout <= 17'h1e0e0;     
      547	:   dout <= 17'h13737;     
      548	:   dout <= 17'h13737;     
      549	:   dout <= 17'h10000;     
      550	:   dout <= 17'h10000;     
      551	:   dout <= 17'h10000;     
      552	:   dout <= 17'h10000;     
      553	:   dout <= 17'h10000;     
      554	:   dout <= 17'h10000;     
      555	:   dout <= 17'h10000;     
      556	:   dout <= 17'h10000;     
      557	:   dout <= 17'h10000;     
      558	:   dout <= 17'h10000;     
      559	:   dout <= 17'h10000;     
      560	:   dout <= 17'h10000;     
      561	:   dout <= 17'h10000;     
      562	:   dout <= 17'h10000;     
      563	:   dout <= 17'h10000;     
      564	:   dout <= 17'h10000;     
      565	:   dout <= 17'h10000;     
      566	:   dout <= 17'h10000;     
      567	:   dout <= 17'h10000;     
      568	:   dout <= 17'h10000;     
      569	:   dout <= 17'h10000;     
      570	:   dout <= 17'h10000;     
      571	:   dout <= 17'h00000;     
      572	:   dout <= 17'h00000;     
      573	:   dout <= 17'h00000;     
      574	:   dout <= 17'h00000;     
      575	:   dout <= 17'h00000;     
      576	:   dout <= 17'h00000;     
      577	:   dout <= 17'h00000;     
      578	:   dout <= 17'h00000;     
      579	:   dout <= 17'h00000;     
      580	:   dout <= 17'h00000;     
      581	:   dout <= 17'h00000;     
      582	:   dout <= 17'h00000;     
      583	:   dout <= 17'h00000;     
      584	:   dout <= 17'h00000;     
      585	:   dout <= 17'h00000;     
      586	:   dout <= 17'h00000;     
      587	:   dout <= 17'h00000;     
      588	:   dout <= 17'h00000;     
      589	:   dout <= 17'h00000;     
      590	:   dout <= 17'h00000;     
      591	:   dout <= 17'h00000;     
      592	:   dout <= 17'h00000;     
      593	:   dout <= 17'h00000;     
      594	:   dout <= 17'h00000;     
      595	:   dout <= 17'h00000;     
      596	:   dout <= 17'h00000;     
      597	:   dout <= 17'h00000;     
      598	:   dout <= 17'h00000;     
      599	:   dout <= 17'h00000;     
      600	:   dout <= 17'h00000;     
      601	:   dout <= 17'h00000;     
      602	:   dout <= 17'h00000;     
      603	:   dout <= 17'h00000;     
      604	:   dout <= 17'h00000;     
      605	:   dout <= 17'h00000;     
      606	:   dout <= 17'h00000;     
      607	:   dout <= 17'h00000;     
      608	:   dout <= 17'h00000;     
      609	:   dout <= 17'h00000;     
      610	:   dout <= 17'h00000;     
      611	:   dout <= 17'h00000;     
      612	:   dout <= 17'h00000;     
      613	:   dout <= 17'h00000;     
      614	:   dout <= 17'h00000;     
      615	:   dout <= 17'h00000;     
      616	:   dout <= 17'h00000;     
      617	:   dout <= 17'h00000;     
      618	:   dout <= 17'h00000;     
      619	:   dout <= 17'h00000;     
      620	:   dout <= 17'h00000;     
      621	:   dout <= 17'h00000;     
      622	:   dout <= 17'h00000;     
      623	:   dout <= 17'h00000;     
      624	:   dout <= 17'h00000;     
      625	:   dout <= 17'h00000;     
      626	:   dout <= 17'h00000;     
      627	:   dout <= 17'h00000;     
      628	:   dout <= 17'h00000;     
      629	:   dout <= 17'h00000;     
      630	:   dout <= 17'h00000;     
      631	:   dout <= 17'h00000;     
      632	:   dout <= 17'h00000;     
      633	:   dout <= 17'h00000;     
      634	:   dout <= 17'h00000;     
      635	:   dout <= 17'h00000;     
      636	:   dout <= 17'h00000;     
      637	:   dout <= 17'h00000;     
      638	:   dout <= 17'h00000;     
      639	:   dout <= 17'h00000;     
      640	:   dout <= 17'h00000;     
      641	:   dout <= 17'h00000;     
      642	:   dout <= 17'h00000;     
      643	:   dout <= 17'h00000;     
      644	:   dout <= 17'h00000;     
      645	:   dout <= 17'h00000;     
      646	:   dout <= 17'h00000;     
      647	:   dout <= 17'h00000;     
      648	:   dout <= 17'h00000;     
      649	:   dout <= 17'h00000;     
      650	:   dout <= 17'h00000;     
      651	:   dout <= 17'h00000;     
      652	:   dout <= 17'h00000;     
      653	:   dout <= 17'h00000;     
      654	:   dout <= 17'h00000;     
      655	:   dout <= 17'h00000;     
      656	:   dout <= 17'h00000;     
      657	:   dout <= 17'h00000;     
      658	:   dout <= 17'h00000;     
      659	:   dout <= 17'h00000;     
      660	:   dout <= 17'h00000;     
      661	:   dout <= 17'h00000;     
      662	:   dout <= 17'h00000;     
      663	:   dout <= 17'h00000;     
      664	:   dout <= 17'h00000;     
      665	:   dout <= 17'h00000;     
      666	:   dout <= 17'h00000;     
      667	:   dout <= 17'h00000;     
      668	:   dout <= 17'h00000;     
      669	:   dout <= 17'h00000;     
      670	:   dout <= 17'h00000;     
      671	:   dout <= 17'h00000;     
      672	:   dout <= 17'h00000;     
      673	:   dout <= 17'h00000;     
      674	:   dout <= 17'h00000;     
      675	:   dout <= 17'h00000;     
      676	:   dout <= 17'h00000;     
      677	:   dout <= 17'h00000;     
      678	:   dout <= 17'h00000;     
      679	:   dout <= 17'h00000;     
      680	:   dout <= 17'h00000;     
      681	:   dout <= 17'h00000;     
      682	:   dout <= 17'h00000;     
      683	:   dout <= 17'h00000;     
      684	:   dout <= 17'h00000;     
      685	:   dout <= 17'h00000;     
      686	:   dout <= 17'h00000;     
      687	:   dout <= 17'h00000;     
      688	:   dout <= 17'h00000;     
      689	:   dout <= 17'h00000;     
      690	:   dout <= 17'h00000;     
      691	:   dout <= 17'h00000;     
      692	:   dout <= 17'h00000;     
      693	:   dout <= 17'h00000;     
      694	:   dout <= 17'h00000;     
      695	:   dout <= 17'h00000;     
      696	:   dout <= 17'h00000;     
      697	:   dout <= 17'h00000;     
      698	:   dout <= 17'h00000;     
      699	:   dout <= 17'h00000;     
      700	:   dout <= 17'h00000;     
      701	:   dout <= 17'h00000;     
      702	:   dout <= 17'h00000;     
      703	:   dout <= 17'h00000;     
      704	:   dout <= 17'h00000;     
      705	:   dout <= 17'h00000;     
      706	:   dout <= 17'h00000;     
      707	:   dout <= 17'h00000;     
      708	:   dout <= 17'h00000;     
      709	:   dout <= 17'h00000;     
      710	:   dout <= 17'h00000;     
      711	:   dout <= 17'h00000;     
      712	:   dout <= 17'h00000;     
      713	:   dout <= 17'h00000;     
      714	:   dout <= 17'h00000;     
      715	:   dout <= 17'h00000;     
      716	:   dout <= 17'h00000;     
      717	:   dout <= 17'h00000;     
      718	:   dout <= 17'h00000;     
      719	:   dout <= 17'h00000;     
      720	:   dout <= 17'h00000;     
      721	:   dout <= 17'h00000;     
      722	:   dout <= 17'h00000;     
      723	:   dout <= 17'h00000;     
      724	:   dout <= 17'h00000;     
      725	:   dout <= 17'h00000;     
      726	:   dout <= 17'h00000;     
      727	:   dout <= 17'h00000;     
      728	:   dout <= 17'h00000;     
      729	:   dout <= 17'h00000;     
      730	:   dout <= 17'h00000;     
      731	:   dout <= 17'h00000;     
      732	:   dout <= 17'h00000;     
      733	:   dout <= 17'h00000;     
      734	:   dout <= 17'h00000;     
      735	:   dout <= 17'h00000;     
      736	:   dout <= 17'h00000;     
      737	:   dout <= 17'h00000;     
      738	:   dout <= 17'h00000;     
      739	:   dout <= 17'h00000;     
      740	:   dout <= 17'h00000;     
      741	:   dout <= 17'h00000;     
      742	:   dout <= 17'h00000;     
      743	:   dout <= 17'h00000;     
      744	:   dout <= 17'h00000;     
      745	:   dout <= 17'h00000;     
      746	:   dout <= 17'h00000;     
      747	:   dout <= 17'h00000;     
      748	:   dout <= 17'h00000;     
      749	:   dout <= 17'h00000;     
      750	:   dout <= 17'h00000;     
      751	:   dout <= 17'h00000;     
      752	:   dout <= 17'h00000;     
      753	:   dout <= 17'h00000;     
      754	:   dout <= 17'h00000;     
      755	:   dout <= 17'h00000;     
      756	:   dout <= 17'h00000;     
      757	:   dout <= 17'h00000;     
      758	:   dout <= 17'h00000;     
      759	:   dout <= 17'h00000;     
      760	:   dout <= 17'h00000;     
      761	:   dout <= 17'h00000;     
      762	:   dout <= 17'h00000;     
      763	:   dout <= 17'h00000;     
      764	:   dout <= 17'h00000;     
      765	:   dout <= 17'h00000;     
      766	:   dout <= 17'h00000;     
      767	:   dout <= 17'h00000;     
      768	:   dout <= 17'h00000;     
      769	:   dout <= 17'h00000;     
      770	:   dout <= 17'h00000;     
      771	:   dout <= 17'h00000;     
      772	:   dout <= 17'h00000;     
      773	:   dout <= 17'h00000;     
      774	:   dout <= 17'h00000;     
      775	:   dout <= 17'h00000;     
      776	:   dout <= 17'h00000;     
      777	:   dout <= 17'h00000;     
      778	:   dout <= 17'h00000;     
      779	:   dout <= 17'h00000;     
      780	:   dout <= 17'h00000;     
      781	:   dout <= 17'h00000;     
      782	:   dout <= 17'h00000;     
      783	:   dout <= 17'h00000;     
      784	:   dout <= 17'h00000;     
      785	:   dout <= 17'h00000;     
      786	:   dout <= 17'h00000;     
      787	:   dout <= 17'h00000;     
      788	:   dout <= 17'h00000;     
      789	:   dout <= 17'h00000;     
      790	:   dout <= 17'h00000;     
      791	:   dout <= 17'h00000;     
      792	:   dout <= 17'h00000;     
      793	:   dout <= 17'h00000;     
      794	:   dout <= 17'h00000;     
      795	:   dout <= 17'h00000;     
      796	:   dout <= 17'h00000;     
      797	:   dout <= 17'h00000;     
      798	:   dout <= 17'h00000;     
      799	:   dout <= 17'h00000;     
      800	:   dout <= 17'h00000;     
      801	:   dout <= 17'h00000;     
      802	:   dout <= 17'h00000;     
      803	:   dout <= 17'h00000;     
      804	:   dout <= 17'h00000;     
      805	:   dout <= 17'h00000;     
      806	:   dout <= 17'h00000;     
      807	:   dout <= 17'h00000;     
      808	:   dout <= 17'h00000;     
      809	:   dout <= 17'h00000;     
      810	:   dout <= 17'h00000;     
      811	:   dout <= 17'h00000;     
      812	:   dout <= 17'h00000;     
      813	:   dout <= 17'h00000;     
      814	:   dout <= 17'h00000;     
      815	:   dout <= 17'h00000;     
      816	:   dout <= 17'h00000;     
      817	:   dout <= 17'h00000;     
      818	:   dout <= 17'h00000;     
      819	:   dout <= 17'h00000;     
      820	:   dout <= 17'h00000;     
      821	:   dout <= 17'h00000;     
      822	:   dout <= 17'h00000;     
      823	:   dout <= 17'h00000;     
      824	:   dout <= 17'h00000;     
      825	:   dout <= 17'h00000;     
      826	:   dout <= 17'h00000;     
      827	:   dout <= 17'h00000;     
      828	:   dout <= 17'h00000;     
      829	:   dout <= 17'h00000;     
      830	:   dout <= 17'h00000;     
      831	:   dout <= 17'h00000;     
      832	:   dout <= 17'h00000;     
      833	:   dout <= 17'h00000;     
      834	:   dout <= 17'h00000;     
      835	:   dout <= 17'h00000;     
      836	:   dout <= 17'h00000;     
      837	:   dout <= 17'h00000;     
      838	:   dout <= 17'h00000;     
      839	:   dout <= 17'h00000;     
      840	:   dout <= 17'h00000;     
      841	:   dout <= 17'h00000;     
      842	:   dout <= 17'h00000;     
      843	:   dout <= 17'h00000;     
      844	:   dout <= 17'h00000;     
      845	:   dout <= 17'h00000;     
      846	:   dout <= 17'h00000;     
      847	:   dout <= 17'h00000;     
      848	:   dout <= 17'h00000;     
      849	:   dout <= 17'h00000;     
      850	:   dout <= 17'h00000;     
      851	:   dout <= 17'h00000;     
      852	:   dout <= 17'h00000;     
      853	:   dout <= 17'h00000;     
      854	:   dout <= 17'h00000;     
      855	:   dout <= 17'h00000;     
      856	:   dout <= 17'h00000;     
      857	:   dout <= 17'h00000;     
      858	:   dout <= 17'h00000;     
      859	:   dout <= 17'h00000;     
      860	:   dout <= 17'h00000;     
      861	:   dout <= 17'h00000;     
      862	:   dout <= 17'h00000;     
      863	:   dout <= 17'h00000;     
      864	:   dout <= 17'h00000;     
      865	:   dout <= 17'h00000;     
      866	:   dout <= 17'h00000;     
      867	:   dout <= 17'h00000;     
      868	:   dout <= 17'h00000;     
      869	:   dout <= 17'h00000;     
      870	:   dout <= 17'h00000;     
      871	:   dout <= 17'h00000;     
      872	:   dout <= 17'h00000;     
      873	:   dout <= 17'h00000;     
      874	:   dout <= 17'h00000;     
      875	:   dout <= 17'h00000;     
      876	:   dout <= 17'h00000;     
      877	:   dout <= 17'h00000;     
      878	:   dout <= 17'h00000;     
      879	:   dout <= 17'h00000;     
      880	:   dout <= 17'h00000;     
      881	:   dout <= 17'h00000;     
      882	:   dout <= 17'h00000;     
      883	:   dout <= 17'h00000;     
      884	:   dout <= 17'h00000;     
      885	:   dout <= 17'h00000;     
      886	:   dout <= 17'h00000;     
      887	:   dout <= 17'h00000;     
      888	:   dout <= 17'h00000;     
      889	:   dout <= 17'h00000;     
      890	:   dout <= 17'h00000;     
      891	:   dout <= 17'h00000;     
      892	:   dout <= 17'h00000;     
      893	:   dout <= 17'h00000;     
      894	:   dout <= 17'h00000;     
      895	:   dout <= 17'h00000;     
      896	:   dout <= 17'h00000;     
      897	:   dout <= 17'h00000;     
      898	:   dout <= 17'h00000;     
      899	:   dout <= 17'h00000;     
      900	:   dout <= 17'h00000;     
      901	:   dout <= 17'h00000;     
      902	:   dout <= 17'h00000;     
      903	:   dout <= 17'h00000;     
      904	:   dout <= 17'h00000;     
      905	:   dout <= 17'h00000;     
      906	:   dout <= 17'h00000;     
      907	:   dout <= 17'h00000;     
      908	:   dout <= 17'h00000;     
      909	:   dout <= 17'h00000;     
      910	:   dout <= 17'h00000;     
      911	:   dout <= 17'h00000;     
      912	:   dout <= 17'h00000;     
      913	:   dout <= 17'h00000;     
      914	:   dout <= 17'h00000;     
      915	:   dout <= 17'h00000;     
      916	:   dout <= 17'h00000;     
      917	:   dout <= 17'h00000;     
      918	:   dout <= 17'h00000;     
      919	:   dout <= 17'h00000;     
      920	:   dout <= 17'h00000;     
      921	:   dout <= 17'h00000;     
      922	:   dout <= 17'h00000;     
      923	:   dout <= 17'h00000;     
      924	:   dout <= 17'h00000;     
      925	:   dout <= 17'h00000;     
      926	:   dout <= 17'h00000;     
      927	:   dout <= 17'h00000;     
      928	:   dout <= 17'h00000;     
      929	:   dout <= 17'h00000;     
      930	:   dout <= 17'h00000;     
      931	:   dout <= 17'h00000;     
      932	:   dout <= 17'h00000;     
      933	:   dout <= 17'h00000;     
      934	:   dout <= 17'h00000;     
      935	:   dout <= 17'h00000;     
      936	:   dout <= 17'h00000;     
      937	:   dout <= 17'h00000;     
      938	:   dout <= 17'h00000;     
      939	:   dout <= 17'h00000;     
      940	:   dout <= 17'h00000;     
      941	:   dout <= 17'h00000;     
      942	:   dout <= 17'h00000;     
      943	:   dout <= 17'h00000;     
      944	:   dout <= 17'h00000;     
      945	:   dout <= 17'h00000;     
      946	:   dout <= 17'h00000;     
      947	:   dout <= 17'h00000;     
      948	:   dout <= 17'h00000;     
      949	:   dout <= 17'h00000;     
      950	:   dout <= 17'h00000;     
      951	:   dout <= 17'h00000;     
      952	:   dout <= 17'h00000;     
      953	:   dout <= 17'h00000;     
      954	:   dout <= 17'h00000;     
      955	:   dout <= 17'h00000;     
      956	:   dout <= 17'h00000;     
      957	:   dout <= 17'h00000;     
      958	:   dout <= 17'h00000;     
      959	:   dout <= 17'h00000;     
      960	:   dout <= 17'h00000;     
      961	:   dout <= 17'h00000;     
      962	:   dout <= 17'h00000;     
      963	:   dout <= 17'h00000;     
      964	:   dout <= 17'h00000;     
      965	:   dout <= 17'h00000;     
      966	:   dout <= 17'h00000;     
      967	:   dout <= 17'h00000;     
      968	:   dout <= 17'h00000;     
      969	:   dout <= 17'h00000;     
      970	:   dout <= 17'h00000;     
      971	:   dout <= 17'h00000;     
      972	:   dout <= 17'h00000;     
      973	:   dout <= 17'h00000;     
      974	:   dout <= 17'h00000;     
      975	:   dout <= 17'h00000;     
      976	:   dout <= 17'h00000;     
      977	:   dout <= 17'h00000;     
      978	:   dout <= 17'h00000;     
      979	:   dout <= 17'h00000;     
      980	:   dout <= 17'h00000;     
      981	:   dout <= 17'h00000;     
      982	:   dout <= 17'h00000;     
      983	:   dout <= 17'h00000;     
      984	:   dout <= 17'h00000;     
      985	:   dout <= 17'h00000;     
      986	:   dout <= 17'h00000;     
      987	:   dout <= 17'h00000;     
      988	:   dout <= 17'h00000;     
      989	:   dout <= 17'h00000;     
      990	:   dout <= 17'h00000;     
      991	:   dout <= 17'h00000;     
      992	:   dout <= 17'h00000;     
      993	:   dout <= 17'h00000;     
      994	:   dout <= 17'h00000;     
      995	:   dout <= 17'h00000;     
      996	:   dout <= 17'h00000;     
      997	:   dout <= 17'h00000;     
      998	:   dout <= 17'h00000;     
      999	:   dout <= 17'h00000;     
      1000	: dout <= 17'h00000;     
      1001	: dout <= 17'h00000;     
      1002	: dout <= 17'h00000;     
      1003	: dout <= 17'h00000;     
      1004	: dout <= 17'h00000;     
      1005	: dout <= 17'h00000;     
      1006	: dout <= 17'h00000;     
      1007	: dout <= 17'h00000;     
      1008	: dout <= 17'h00000;     
      1009	: dout <= 17'h00000;     
      1010	: dout <= 17'h00000;     
      1011	: dout <= 17'h00000;     
      1012	: dout <= 17'h00000;     
      1013	: dout <= 17'h00000;     
      1014	: dout <= 17'h00000;     
      1015	: dout <= 17'h00000;     
      1016	: dout <= 17'h00000;     
      1017	: dout <= 17'h00000;     
      1018	: dout <= 17'h00000;     
      1019	: dout <= 17'h00000;     
      1020	: dout <= 17'h00000;     
      1021	: dout <= 17'h00000;     
      1022	: dout <= 17'h00000;     
      default:dout <= 17'h00000;
    endcase
  end
endmodule

